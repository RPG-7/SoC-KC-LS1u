module alu74181(a,b,cin, s,m, f, cout, eqv, g,p);


input [3:0] a,b,s;
input cin;
input m;
output [3:0] f;
output g , p;
output cout, eqv;   

wire	SYNTHESIZED_WIRE_117;
wire	SYNTHESIZED_WIRE_118;
wire	SYNTHESIZED_WIRE_119;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_128;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_98;
wire	SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_101;
wire	SYNTHESIZED_WIRE_102;
wire	SYNTHESIZED_WIRE_103;
wire	SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_116;
wire	SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_112;
wire	SYNTHESIZED_WIRE_113;
wire	SYNTHESIZED_WIRE_114;
wire	SYNTHESIZED_WIRE_115;

assign	f[1] = SYNTHESIZED_WIRE_113;
assign	f[2] = SYNTHESIZED_WIRE_112;
assign	f[3] = SYNTHESIZED_WIRE_111;
assign	g = SYNTHESIZED_WIRE_96;
assign	f[0] = SYNTHESIZED_WIRE_114;

assign	SYNTHESIZED_WIRE_14 = s[0] & b[1];

assign	SYNTHESIZED_WIRE_15 = SYNTHESIZED_WIRE_117 & s[1];

assign	SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_117 & s[2] & a[1];

assign	SYNTHESIZED_WIRE_20 = a[1] & s[3] & b[1];

assign	SYNTHESIZED_WIRE_16 = s[0] & b[2];

assign	SYNTHESIZED_WIRE_17 = SYNTHESIZED_WIRE_118 & s[1];

assign	SYNTHESIZED_WIRE_23 = SYNTHESIZED_WIRE_118 & s[2] & a[2];

assign	SYNTHESIZED_WIRE_22 = a[2] & s[3] & b[2];

assign	SYNTHESIZED_WIRE_26 = s[0] & b[3];

assign	SYNTHESIZED_WIRE_27 = SYNTHESIZED_WIRE_119 & s[1];

assign	SYNTHESIZED_WIRE_29 = SYNTHESIZED_WIRE_119 & s[2] & a[3];

assign	SYNTHESIZED_WIRE_28 = a[3] & s[3] & b[3];

assign	SYNTHESIZED_WIRE_119 =  ~b[3];

assign	SYNTHESIZED_WIRE_129 =  ~b[0];

assign	SYNTHESIZED_WIRE_117 =  ~b[1];

assign	SYNTHESIZED_WIRE_118 =  ~b[2];

assign	SYNTHESIZED_WIRE_6 = ~(a[0] | SYNTHESIZED_WIRE_12 | SYNTHESIZED_WIRE_13);

assign	SYNTHESIZED_WIRE_8 = ~(a[1] | SYNTHESIZED_WIRE_14 | SYNTHESIZED_WIRE_15);

assign	SYNTHESIZED_WIRE_10 = ~(a[2] | SYNTHESIZED_WIRE_16 | SYNTHESIZED_WIRE_17);

assign	SYNTHESIZED_WIRE_7 = ~(SYNTHESIZED_WIRE_18 | SYNTHESIZED_WIRE_19);

assign	SYNTHESIZED_WIRE_9 = ~(SYNTHESIZED_WIRE_20 | SYNTHESIZED_WIRE_21);

assign	SYNTHESIZED_WIRE_11 = ~(SYNTHESIZED_WIRE_22 | SYNTHESIZED_WIRE_23);

assign	SYNTHESIZED_WIRE_25 = ~(a[3] | SYNTHESIZED_WIRE_26 | SYNTHESIZED_WIRE_27);

assign	SYNTHESIZED_WIRE_24 = ~(SYNTHESIZED_WIRE_28 | SYNTHESIZED_WIRE_29);

assign	SYNTHESIZED_WIRE_101 = SYNTHESIZED_WIRE_7 ^ SYNTHESIZED_WIRE_6;

assign	SYNTHESIZED_WIRE_103 = SYNTHESIZED_WIRE_9 ^ SYNTHESIZED_WIRE_8;

assign	SYNTHESIZED_WIRE_105 = SYNTHESIZED_WIRE_11 ^ SYNTHESIZED_WIRE_10;

assign	SYNTHESIZED_WIRE_94 = SYNTHESIZED_WIRE_24 ^ SYNTHESIZED_WIRE_25;

assign	SYNTHESIZED_WIRE_56 = SYNTHESIZED_WIRE_24 & SYNTHESIZED_WIRE_10;

assign	SYNTHESIZED_WIRE_57 = SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_24;

assign	SYNTHESIZED_WIRE_12 = s[0] & b[0];

assign	p = ~(SYNTHESIZED_WIRE_24 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_7);

assign	SYNTHESIZED_WIRE_97 = ~(SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_24 & cin & cin);

assign	SYNTHESIZED_WIRE_58 = SYNTHESIZED_WIRE_24 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_6;

assign	SYNTHESIZED_WIRE_96 = ~(SYNTHESIZED_WIRE_25 | SYNTHESIZED_WIRE_56 | SYNTHESIZED_WIRE_57 | SYNTHESIZED_WIRE_58);

assign	SYNTHESIZED_WIRE_102 = ~(cin & SYNTHESIZED_WIRE_128);

assign	SYNTHESIZED_WIRE_99 = SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_98 = SYNTHESIZED_WIRE_128 & SYNTHESIZED_WIRE_7 & cin;

assign	SYNTHESIZED_WIRE_90 = SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_91 = SYNTHESIZED_WIRE_128 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_9;

assign	SYNTHESIZED_WIRE_92 = cin & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_13 = SYNTHESIZED_WIRE_129 & s[1];

assign	SYNTHESIZED_WIRE_89 = SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_88 = SYNTHESIZED_WIRE_128 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_11;

assign	SYNTHESIZED_WIRE_87 = SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_86 = cin & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_9 & cin & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_93 = ~(SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_88 | SYNTHESIZED_WIRE_89);

assign	SYNTHESIZED_WIRE_116 = ~(SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_92);

assign	SYNTHESIZED_WIRE_111 = SYNTHESIZED_WIRE_94 ^ SYNTHESIZED_WIRE_93;

assign	cout = ~(SYNTHESIZED_WIRE_96 & SYNTHESIZED_WIRE_97);

assign	SYNTHESIZED_WIRE_115 = ~(SYNTHESIZED_WIRE_98 | SYNTHESIZED_WIRE_99);

assign	SYNTHESIZED_WIRE_19 = SYNTHESIZED_WIRE_129 & s[2] & a[0];

assign	SYNTHESIZED_WIRE_114 = SYNTHESIZED_WIRE_101 ^ SYNTHESIZED_WIRE_102;

assign	SYNTHESIZED_WIRE_113 = SYNTHESIZED_WIRE_103 ^ SYNTHESIZED_WIRE_115;

assign	SYNTHESIZED_WIRE_112 = SYNTHESIZED_WIRE_105 ^ SYNTHESIZED_WIRE_116;

assign	eqv = SYNTHESIZED_WIRE_111 & SYNTHESIZED_WIRE_112 & SYNTHESIZED_WIRE_113 & SYNTHESIZED_WIRE_114;

assign	SYNTHESIZED_WIRE_18 = a[0] & s[3] & b[0];

assign	SYNTHESIZED_WIRE_128 =  ~m;
endmodule
