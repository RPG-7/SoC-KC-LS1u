module cdma
(
    
);



endmodule
