module hbus_mux
(

);


endmodule
