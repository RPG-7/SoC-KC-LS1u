/* Verilog module written by vlog2Verilog (qflow) */

module KC_LS1u(
    input WAIT,
    input clk,
    output [23:0] daddr,
    input [7:0] ddata_i,
    output [7:0] ddata_o,
    output dwrite,
    output [23:0] iaddr,
    input [15:0] instr,
    input rst
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire [7:0] C ;
wire [7:0] D ;
wire _588_ ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _19_ ;
wire _512_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _415_ ;
wire _95_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _262_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _259_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_121  ;
wire _488_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_108  ;
wire _412_ ;
wire _92_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _197_ ;
wire _7_ ;
wire WAIT ;
wire _503_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _215_ ;
wire _444_ ;
wire _253_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_10  ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_109  ;
wire _212_ ;
wire _441_ ;
wire _250_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire _285_ ;
wire _1_ ;
wire [3:0] \ALU_H4.b  ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_106  ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _206_ ;
wire _435_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _432_ ;
wire _241_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _93__bF$buf0 ;
wire _93__bF$buf1 ;
wire _93__bF$buf2 ;
wire _93__bF$buf3 ;
wire _93__bF$buf4 ;
wire _429_ ;
wire _182_ ;
wire _238_ ;
wire _467_ ;
wire _276_ ;
wire _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire _523_ ;
wire _103_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _370_ ;
wire _426_ ;
wire _235_ ;
wire _464_ ;
wire WAIT_bF$buf0 ;
wire WAIT_bF$buf1 ;
wire WAIT_bF$buf2 ;
wire WAIT_bF$buf3 ;
wire WAIT_bF$buf4 ;
wire _273_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire [15:0] instr ;
wire _30_ ;
wire _367_ ;
wire _176_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_122  ;
wire _499_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _423_ ;
wire _232_ ;
wire _461_ ;
wire _517_ ;
wire _270_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _173_ ;
wire _229_ ;
wire _458_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _420_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_126  ;
wire _514_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire [7:0] _590_ ;
wire _170_ ;
wire _226_ ;
wire _455_ ;
wire _264_ ;
wire \ALU_H4.p  ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire [3:0] \ALU_L4.b  ;
wire \ALU_L4.SYNTHESIZED_WIRE_123  ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _320_ ;
wire _56_ ;
wire _414_ ;
wire _94_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _261_ ;
wire _317_ ;
wire _490_ ;
wire [7:0] ddata_i ;
wire [7:0] ddata_o ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_93  ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_110  ;
wire _258_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_120  ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire \ALU_H4.eqv  ;
wire _53_ ;
wire _199_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_107  ;
wire _411_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_104  ;
wire \ALU_L4.SYNTHESIZED_WIRE_11  ;
wire _6_ ;
wire _502_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _214_ ;
wire _443_ ;
wire _252_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire rst ;
wire _290_ ;
wire _346_ ;
wire _351__bF$buf0 ;
wire _351__bF$buf1 ;
wire _351__bF$buf2 ;
wire _351__bF$buf3 ;
wire _351__bF$buf4 ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_108  ;
wire _211_ ;
wire _440_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire [3:0] \ALU_H4.a  ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _205_ ;
wire _434_ ;
wire _243_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_127  ;
wire _431_ ;
wire _240_ ;
wire _525_ ;
wire _105_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _237_ ;
wire _466_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire [23:0] iaddr ;
wire _425_ ;
wire [23:0] daddr ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _272_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _175_ ;
wire dwrite ;
wire \ALU_H4.SYNTHESIZED_WIRE_121  ;
wire _269_ ;
wire \ALU_H4.cout  ;
wire _498_ ;
wire _26_ ;
wire _64_ ;
wire _422_ ;
wire _231_ ;
wire _460_ ;
wire _516_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire [23:0] _592_ ;
wire _172_ ;
wire _228_ ;
wire _457_ ;
wire _266_ ;
wire _495_ ;
wire _161__bF$buf0 ;
wire _161__bF$buf1 ;
wire _161__bF$buf2 ;
wire _161__bF$buf3 ;
wire _161__bF$buf4 ;
wire _161__bF$buf5 ;
wire _161__bF$buf6 ;
wire _161__bF$buf7 ;
wire _23_ ;
wire [23:0] _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _513_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire _225_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_96  ;
wire _454_ ;
wire _263_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire [3:0] \ALU_L4.a  ;
wire \ALU_L4.SYNTHESIZED_WIRE_122  ;
wire _489_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_109  ;
wire _413_ ;
wire _93_ ;
wire _222_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_93  ;
wire _451_ ;
wire _507_ ;
wire _260_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _198_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_106  ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _216_ ;
wire _445_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_11  ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_10  ;
wire _5_ ;
wire _501_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _213_ ;
wire _442_ ;
wire _251_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _248_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_110  ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_107  ;
wire _210_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_104  ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _204_ ;
wire _433_ ;
wire _242_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _239_ ;
wire _468_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_126  ;
wire _430_ ;
wire _524_ ;
wire _104_ ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _236_ ;
wire _465_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _177_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_123  ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _330_ ;
wire _66_ ;
wire _424_ ;
wire _233_ ;
wire _462_ ;
wire _518_ ;
wire _271_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _174_ ;
wire \ALU_L4.eqv  ;
wire _459_ ;
wire \ALU_H4.SYNTHESIZED_WIRE_120  ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _63_ ;
wire _421_ ;
wire \ALU_L4.SYNTHESIZED_WIRE_127  ;
wire _230_ ;
wire _515_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _227_ ;
wire _456_ ;
wire _265_ ;
wire _494_ ;
wire _0__bF$buf0 ;
wire _0__bF$buf1 ;
wire _0__bF$buf2 ;
wire _0__bF$buf3 ;
wire _22_ ;
wire _359_ ;

BUFX2 BUFX2_insert35 (
    .A(_351_),
    .Y(_351__bF$buf0)
);

BUFX2 BUFX2_insert34 (
    .A(_351_),
    .Y(_351__bF$buf1)
);

BUFX2 BUFX2_insert33 (
    .A(_351_),
    .Y(_351__bF$buf2)
);

BUFX2 BUFX2_insert32 (
    .A(_351_),
    .Y(_351__bF$buf3)
);

BUFX2 BUFX2_insert31 (
    .A(_351_),
    .Y(_351__bF$buf4)
);

BUFX2 BUFX2_insert30 (
    .A(_93_),
    .Y(_93__bF$buf0)
);

BUFX2 BUFX2_insert29 (
    .A(_93_),
    .Y(_93__bF$buf1)
);

BUFX2 BUFX2_insert28 (
    .A(_93_),
    .Y(_93__bF$buf2)
);

BUFX2 BUFX2_insert27 (
    .A(_93_),
    .Y(_93__bF$buf3)
);

BUFX2 BUFX2_insert26 (
    .A(_93_),
    .Y(_93__bF$buf4)
);

BUFX2 BUFX2_insert25 (
    .A(_0_),
    .Y(_0__bF$buf0)
);

BUFX2 BUFX2_insert24 (
    .A(_0_),
    .Y(_0__bF$buf1)
);

BUFX2 BUFX2_insert23 (
    .A(_0_),
    .Y(_0__bF$buf2)
);

BUFX2 BUFX2_insert22 (
    .A(_0_),
    .Y(_0__bF$buf3)
);

BUFX2 BUFX2_insert21 (
    .A(_161_),
    .Y(_161__bF$buf0)
);

BUFX2 BUFX2_insert20 (
    .A(_161_),
    .Y(_161__bF$buf1)
);

BUFX2 BUFX2_insert19 (
    .A(_161_),
    .Y(_161__bF$buf2)
);

BUFX2 BUFX2_insert18 (
    .A(_161_),
    .Y(_161__bF$buf3)
);

BUFX2 BUFX2_insert17 (
    .A(_161_),
    .Y(_161__bF$buf4)
);

BUFX2 BUFX2_insert16 (
    .A(_161_),
    .Y(_161__bF$buf5)
);

BUFX2 BUFX2_insert15 (
    .A(_161_),
    .Y(_161__bF$buf6)
);

BUFX2 BUFX2_insert14 (
    .A(_161_),
    .Y(_161__bF$buf7)
);

CLKBUF1 CLKBUF1_insert13 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert11 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert10 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert9 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert8 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert7 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert6 (
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert5 (
    .A(clk),
    .Y(clk_bF$buf8)
);

BUFX2 BUFX2_insert4 (
    .A(WAIT),
    .Y(WAIT_bF$buf0)
);

BUFX2 BUFX2_insert3 (
    .A(WAIT),
    .Y(WAIT_bF$buf1)
);

BUFX2 BUFX2_insert2 (
    .A(WAIT),
    .Y(WAIT_bF$buf2)
);

BUFX2 BUFX2_insert1 (
    .A(WAIT),
    .Y(WAIT_bF$buf3)
);

BUFX2 BUFX2_insert0 (
    .A(WAIT),
    .Y(WAIT_bF$buf4)
);

NAND2X1 _1000_ (
    .A(_368_),
    .B(_420_),
    .Y(_421_)
);

NOR2X1 _1001_ (
    .A(_408_),
    .B(_421_),
    .Y(_422_)
);

NAND2X1 _1002_ (
    .A(_592_[10]),
    .B(_422_),
    .Y(_423_)
);

XNOR2X1 _1003_ (
    .A(_423_),
    .B(_592_[11]),
    .Y(_424_)
);

MUX2X1 _1004_ (
    .A(_424_),
    .B(_589_[11]),
    .S(_351__bF$buf4),
    .Y(_425_)
);

OAI21X1 _1005_ (
    .A(_425_),
    .B(WAIT_bF$buf4),
    .C(_419_),
    .Y(_77_)
);

INVX2 _1006_ (
    .A(_592_[12]),
    .Y(_426_)
);

NAND2X1 _1007_ (
    .A(_592_[10]),
    .B(_592_[11]),
    .Y(_427_)
);

NOR2X1 _1008_ (
    .A(_408_),
    .B(_427_),
    .Y(_428_)
);

INVX1 _1009_ (
    .A(_428_),
    .Y(_429_)
);

OAI21X1 _1010_ (
    .A(_401_),
    .B(_429_),
    .C(_426_),
    .Y(_430_)
);

NAND3X1 _1011_ (
    .A(_592_[12]),
    .B(_428_),
    .C(_395_),
    .Y(_431_)
);

AOI21X1 _1012_ (
    .A(_430_),
    .B(_431_),
    .C(_353_),
    .Y(_432_)
);

OAI21X1 _1013_ (
    .A(_351__bF$buf3),
    .B(_589_[12]),
    .C(_93__bF$buf4),
    .Y(_433_)
);

OAI22X1 _1014_ (
    .A(_93__bF$buf3),
    .B(_426_),
    .C(_432_),
    .D(_433_),
    .Y(_78_)
);

NAND3X1 _1015_ (
    .A(_368_),
    .B(_420_),
    .C(_428_),
    .Y(_434_)
);

OAI21X1 _1016_ (
    .A(_434_),
    .B(_426_),
    .C(_592_[13]),
    .Y(_435_)
);

INVX1 _1017_ (
    .A(_592_[13]),
    .Y(_436_)
);

NOR2X1 _1018_ (
    .A(_426_),
    .B(_434_),
    .Y(_437_)
);

NAND2X1 _1019_ (
    .A(_436_),
    .B(_437_),
    .Y(_438_)
);

NAND3X1 _1020_ (
    .A(_435_),
    .B(_438_),
    .C(_351__bF$buf2),
    .Y(_439_)
);

OAI21X1 _1021_ (
    .A(_589_[13]),
    .B(_351__bF$buf1),
    .C(_439_),
    .Y(_440_)
);

NAND2X1 _1022_ (
    .A(WAIT_bF$buf3),
    .B(_592_[13]),
    .Y(_441_)
);

OAI21X1 _1023_ (
    .A(_440_),
    .B(WAIT_bF$buf2),
    .C(_441_),
    .Y(_79_)
);

INVX2 _1024_ (
    .A(_592_[14]),
    .Y(_442_)
);

NAND2X1 _1025_ (
    .A(_592_[12]),
    .B(_592_[13]),
    .Y(_443_)
);

OR2X2 _1026_ (
    .A(_434_),
    .B(_443_),
    .Y(_444_)
);

NOR2X1 _1027_ (
    .A(_592_[14]),
    .B(_444_),
    .Y(_445_)
);

NOR2X1 _1028_ (
    .A(_443_),
    .B(_434_),
    .Y(_446_)
);

NOR2X1 _1029_ (
    .A(_442_),
    .B(_446_),
    .Y(_447_)
);

NOR2X1 _1030_ (
    .A(_447_),
    .B(_445_),
    .Y(_448_)
);

AND2X2 _1031_ (
    .A(_448_),
    .B(_351__bF$buf0),
    .Y(_449_)
);

OAI21X1 _1032_ (
    .A(_351__bF$buf4),
    .B(_589_[14]),
    .C(_93__bF$buf2),
    .Y(_450_)
);

OAI22X1 _1033_ (
    .A(_93__bF$buf1),
    .B(_442_),
    .C(_449_),
    .D(_450_),
    .Y(_80_)
);

INVX1 _1034_ (
    .A(_592_[15]),
    .Y(_451_)
);

OAI21X1 _1035_ (
    .A(_444_),
    .B(_442_),
    .C(_592_[15]),
    .Y(_452_)
);

NAND3X1 _1036_ (
    .A(_592_[14]),
    .B(_451_),
    .C(_446_),
    .Y(_453_)
);

NAND3X1 _1037_ (
    .A(_452_),
    .B(_453_),
    .C(_389_),
    .Y(_454_)
);

INVX1 _1038_ (
    .A(_589_[15]),
    .Y(_455_)
);

AOI21X1 _1039_ (
    .A(_346_),
    .B(_348_),
    .C(_97_),
    .Y(_456_)
);

NAND3X1 _1040_ (
    .A(_455_),
    .B(_102_),
    .C(_456_),
    .Y(_457_)
);

NAND3X1 _1041_ (
    .A(_93__bF$buf0),
    .B(_457_),
    .C(_454_),
    .Y(_458_)
);

OAI21X1 _1042_ (
    .A(_93__bF$buf4),
    .B(_451_),
    .C(_458_),
    .Y(_81_)
);

NAND2X1 _1043_ (
    .A(_592_[14]),
    .B(_592_[15]),
    .Y(_459_)
);

NOR2X1 _1044_ (
    .A(_443_),
    .B(_459_),
    .Y(_460_)
);

NAND2X1 _1045_ (
    .A(_428_),
    .B(_460_),
    .Y(_461_)
);

NOR2X1 _1046_ (
    .A(_401_),
    .B(_461_),
    .Y(_462_)
);

NOR2X1 _1047_ (
    .A(_592_[16]),
    .B(_462_),
    .Y(_463_)
);

INVX1 _1048_ (
    .A(_592_[16]),
    .Y(_464_)
);

AND2X2 _1049_ (
    .A(_428_),
    .B(_460_),
    .Y(_465_)
);

NAND2X1 _1050_ (
    .A(_465_),
    .B(_395_),
    .Y(_466_)
);

NOR2X1 _1051_ (
    .A(_464_),
    .B(_466_),
    .Y(_467_)
);

OAI21X1 _1052_ (
    .A(_467_),
    .B(_463_),
    .C(_351__bF$buf3),
    .Y(_468_)
);

OAI21X1 _1053_ (
    .A(_589_[16]),
    .B(_351__bF$buf2),
    .C(_468_),
    .Y(_469_)
);

NAND2X1 _1054_ (
    .A(WAIT_bF$buf1),
    .B(_592_[16]),
    .Y(_470_)
);

OAI21X1 _1055_ (
    .A(_469_),
    .B(WAIT_bF$buf0),
    .C(_470_),
    .Y(_82_)
);

NAND2X1 _1056_ (
    .A(_592_[16]),
    .B(_462_),
    .Y(_471_)
);

XNOR2X1 _1057_ (
    .A(_471_),
    .B(_592_[17]),
    .Y(_472_)
);

OR2X2 _1058_ (
    .A(_351__bF$buf1),
    .B(_589_[17]),
    .Y(_473_)
);

OAI21X1 _1059_ (
    .A(_472_),
    .B(_353_),
    .C(_473_),
    .Y(_474_)
);

NAND2X1 _1060_ (
    .A(WAIT_bF$buf4),
    .B(_592_[17]),
    .Y(_475_)
);

OAI21X1 _1061_ (
    .A(_474_),
    .B(WAIT_bF$buf3),
    .C(_475_),
    .Y(_83_)
);

INVX2 _1062_ (
    .A(_592_[18]),
    .Y(_476_)
);

NAND2X1 _1063_ (
    .A(_592_[16]),
    .B(_592_[17]),
    .Y(_477_)
);

OAI21X1 _1064_ (
    .A(_466_),
    .B(_477_),
    .C(_476_),
    .Y(_478_)
);

NOR2X1 _1065_ (
    .A(_477_),
    .B(_466_),
    .Y(_479_)
);

NAND2X1 _1066_ (
    .A(_592_[18]),
    .B(_479_),
    .Y(_480_)
);

AOI21X1 _1067_ (
    .A(_478_),
    .B(_480_),
    .C(_353_),
    .Y(_481_)
);

OAI21X1 _1068_ (
    .A(_351__bF$buf0),
    .B(_589_[18]),
    .C(_93__bF$buf3),
    .Y(_482_)
);

OAI22X1 _1069_ (
    .A(_93__bF$buf2),
    .B(_476_),
    .C(_481_),
    .D(_482_),
    .Y(_84_)
);

INVX1 _1070_ (
    .A(_592_[19]),
    .Y(_483_)
);

AND2X2 _1071_ (
    .A(_368_),
    .B(_420_),
    .Y(_484_)
);

INVX1 _1072_ (
    .A(_477_),
    .Y(_485_)
);

NAND3X1 _1073_ (
    .A(_485_),
    .B(_484_),
    .C(_465_),
    .Y(_486_)
);

OAI21X1 _1074_ (
    .A(_486_),
    .B(_476_),
    .C(_592_[19]),
    .Y(_487_)
);

NOR3X1 _1075_ (
    .A(_421_),
    .B(_477_),
    .C(_461_),
    .Y(_488_)
);

NAND3X1 _1076_ (
    .A(_592_[18]),
    .B(_483_),
    .C(_488_),
    .Y(_489_)
);

NAND3X1 _1077_ (
    .A(_487_),
    .B(_489_),
    .C(_389_),
    .Y(_490_)
);

INVX1 _1078_ (
    .A(_589_[19]),
    .Y(_491_)
);

NAND3X1 _1079_ (
    .A(_491_),
    .B(_102_),
    .C(_456_),
    .Y(_492_)
);

NAND3X1 _1080_ (
    .A(_93__bF$buf1),
    .B(_492_),
    .C(_490_),
    .Y(_493_)
);

OAI21X1 _1081_ (
    .A(_93__bF$buf0),
    .B(_483_),
    .C(_493_),
    .Y(_85_)
);

INVX1 _1082_ (
    .A(_592_[20]),
    .Y(_494_)
);

NAND2X1 _1083_ (
    .A(_592_[18]),
    .B(_592_[19]),
    .Y(_495_)
);

NOR2X1 _1084_ (
    .A(_477_),
    .B(_495_),
    .Y(_496_)
);

INVX1 _1085_ (
    .A(_496_),
    .Y(_497_)
);

OAI21X1 _1086_ (
    .A(_466_),
    .B(_497_),
    .C(_494_),
    .Y(_498_)
);

NOR3X1 _1087_ (
    .A(_461_),
    .B(_497_),
    .C(_407_),
    .Y(_499_)
);

NAND2X1 _1088_ (
    .A(_592_[20]),
    .B(_499_),
    .Y(_500_)
);

AOI21X1 _1089_ (
    .A(_498_),
    .B(_500_),
    .C(_353_),
    .Y(_501_)
);

OAI21X1 _1090_ (
    .A(_351__bF$buf4),
    .B(_589_[20]),
    .C(_93__bF$buf4),
    .Y(_502_)
);

OAI22X1 _1091_ (
    .A(_93__bF$buf3),
    .B(_494_),
    .C(_501_),
    .D(_502_),
    .Y(_86_)
);

INVX1 _1092_ (
    .A(_592_[21]),
    .Y(_503_)
);

NAND3X1 _1093_ (
    .A(_465_),
    .B(_496_),
    .C(_395_),
    .Y(_504_)
);

NAND2X1 _1094_ (
    .A(_592_[20]),
    .B(_592_[21]),
    .Y(_505_)
);

NOR2X1 _1095_ (
    .A(_505_),
    .B(_504_),
    .Y(_506_)
);

AOI21X1 _1096_ (
    .A(_503_),
    .B(_500_),
    .C(_506_),
    .Y(_507_)
);

NOR2X1 _1097_ (
    .A(_353_),
    .B(_507_),
    .Y(_508_)
);

OAI21X1 _1098_ (
    .A(_351__bF$buf3),
    .B(_589_[21]),
    .C(_93__bF$buf2),
    .Y(_509_)
);

OAI22X1 _1099_ (
    .A(_93__bF$buf1),
    .B(_503_),
    .C(_508_),
    .D(_509_),
    .Y(_87_)
);

INVX1 _1100_ (
    .A(_592_[22]),
    .Y(_510_)
);

OAI21X1 _1101_ (
    .A(_504_),
    .B(_505_),
    .C(_510_),
    .Y(_511_)
);

INVX1 _1102_ (
    .A(_505_),
    .Y(_512_)
);

NAND3X1 _1103_ (
    .A(_592_[22]),
    .B(_512_),
    .C(_499_),
    .Y(_513_)
);

AOI21X1 _1104_ (
    .A(_513_),
    .B(_511_),
    .C(_353_),
    .Y(_514_)
);

OAI21X1 _1105_ (
    .A(_351__bF$buf2),
    .B(_589_[22]),
    .C(_93__bF$buf0),
    .Y(_515_)
);

OAI22X1 _1106_ (
    .A(_93__bF$buf4),
    .B(_510_),
    .C(_514_),
    .D(_515_),
    .Y(_88_)
);

NAND2X1 _1107_ (
    .A(WAIT_bF$buf2),
    .B(_592_[23]),
    .Y(_516_)
);

INVX1 _1108_ (
    .A(_592_[23]),
    .Y(_517_)
);

NAND2X1 _1109_ (
    .A(_517_),
    .B(_513_),
    .Y(_518_)
);

NAND3X1 _1110_ (
    .A(_592_[22]),
    .B(_592_[23]),
    .C(_506_),
    .Y(_519_)
);

AOI21X1 _1111_ (
    .A(_518_),
    .B(_519_),
    .C(_353_),
    .Y(_520_)
);

OAI21X1 _1112_ (
    .A(_351__bF$buf1),
    .B(_589_[23]),
    .C(_93__bF$buf3),
    .Y(_521_)
);

OAI21X1 _1113_ (
    .A(_520_),
    .B(_521_),
    .C(_516_),
    .Y(_89_)
);

INVX1 _1114_ (
    .A(_333_),
    .Y(_33_)
);

DFFPOSX1 _1115_ (
    .CLK(clk_bF$buf8),
    .D(_1_),
    .Q(\ALU_L4.a [0])
);

DFFPOSX1 _1116_ (
    .CLK(clk_bF$buf7),
    .D(_2_),
    .Q(\ALU_L4.a [1])
);

DFFPOSX1 _1117_ (
    .CLK(clk_bF$buf6),
    .D(_3_),
    .Q(\ALU_L4.a [2])
);

DFFPOSX1 _1118_ (
    .CLK(clk_bF$buf5),
    .D(_4_),
    .Q(\ALU_L4.a [3])
);

DFFPOSX1 _1119_ (
    .CLK(clk_bF$buf4),
    .D(_5_),
    .Q(\ALU_H4.a [0])
);

DFFPOSX1 _1120_ (
    .CLK(clk_bF$buf3),
    .D(_6_),
    .Q(\ALU_H4.a [1])
);

DFFPOSX1 _1121_ (
    .CLK(clk_bF$buf2),
    .D(_7_),
    .Q(\ALU_H4.a [2])
);

DFFPOSX1 _1122_ (
    .CLK(clk_bF$buf1),
    .D(_8_),
    .Q(\ALU_H4.a [3])
);

DFFPOSX1 _1123_ (
    .CLK(clk_bF$buf0),
    .D(_9_),
    .Q(\ALU_L4.b [0])
);

DFFPOSX1 _1124_ (
    .CLK(clk_bF$buf8),
    .D(_10_),
    .Q(\ALU_L4.b [1])
);

DFFPOSX1 _1125_ (
    .CLK(clk_bF$buf7),
    .D(_11_),
    .Q(\ALU_L4.b [2])
);

DFFPOSX1 _1126_ (
    .CLK(clk_bF$buf6),
    .D(_12_),
    .Q(\ALU_L4.b [3])
);

DFFPOSX1 _1127_ (
    .CLK(clk_bF$buf5),
    .D(_13_),
    .Q(\ALU_H4.b [0])
);

DFFPOSX1 _1128_ (
    .CLK(clk_bF$buf4),
    .D(_14_),
    .Q(\ALU_H4.b [1])
);

DFFPOSX1 _1129_ (
    .CLK(clk_bF$buf3),
    .D(_15_),
    .Q(\ALU_H4.b [2])
);

DFFPOSX1 _1130_ (
    .CLK(clk_bF$buf2),
    .D(_16_),
    .Q(\ALU_H4.b [3])
);

DFFPOSX1 _1131_ (
    .CLK(clk_bF$buf1),
    .D(_17_),
    .Q(C[0])
);

DFFPOSX1 _1132_ (
    .CLK(clk_bF$buf0),
    .D(_18_),
    .Q(C[1])
);

DFFPOSX1 _1133_ (
    .CLK(clk_bF$buf8),
    .D(_19_),
    .Q(C[2])
);

DFFPOSX1 _1134_ (
    .CLK(clk_bF$buf7),
    .D(_20_),
    .Q(C[3])
);

DFFPOSX1 _1135_ (
    .CLK(clk_bF$buf6),
    .D(_21_),
    .Q(C[4])
);

DFFPOSX1 _1136_ (
    .CLK(clk_bF$buf5),
    .D(_22_),
    .Q(C[5])
);

DFFPOSX1 _1137_ (
    .CLK(clk_bF$buf4),
    .D(_23_),
    .Q(C[6])
);

DFFPOSX1 _1138_ (
    .CLK(clk_bF$buf3),
    .D(_24_),
    .Q(C[7])
);

DFFPOSX1 _1139_ (
    .CLK(clk_bF$buf2),
    .D(_25_),
    .Q(D[0])
);

DFFPOSX1 _1140_ (
    .CLK(clk_bF$buf1),
    .D(_26_),
    .Q(D[1])
);

DFFPOSX1 _1141_ (
    .CLK(clk_bF$buf0),
    .D(_27_),
    .Q(D[2])
);

DFFPOSX1 _1142_ (
    .CLK(clk_bF$buf8),
    .D(_28_),
    .Q(D[3])
);

DFFPOSX1 _1143_ (
    .CLK(clk_bF$buf7),
    .D(_29_),
    .Q(D[4])
);

DFFPOSX1 _1144_ (
    .CLK(clk_bF$buf6),
    .D(_30_),
    .Q(D[5])
);

DFFPOSX1 _1145_ (
    .CLK(clk_bF$buf5),
    .D(_31_),
    .Q(D[6])
);

DFFPOSX1 _1146_ (
    .CLK(clk_bF$buf4),
    .D(_32_),
    .Q(D[7])
);

DFFPOSX1 _1147_ (
    .CLK(clk_bF$buf3),
    .D(_33_),
    .Q(_591_)
);

DFFPOSX1 _1148_ (
    .CLK(clk_bF$buf2),
    .D(_34_),
    .Q(_589_[0])
);

DFFPOSX1 _1149_ (
    .CLK(clk_bF$buf1),
    .D(_35_),
    .Q(_589_[1])
);

DFFPOSX1 _1150_ (
    .CLK(clk_bF$buf0),
    .D(_36_),
    .Q(_589_[2])
);

DFFPOSX1 _1151_ (
    .CLK(clk_bF$buf8),
    .D(_37_),
    .Q(_589_[3])
);

DFFPOSX1 _1152_ (
    .CLK(clk_bF$buf7),
    .D(_38_),
    .Q(_589_[4])
);

DFFPOSX1 _1153_ (
    .CLK(clk_bF$buf6),
    .D(_39_),
    .Q(_589_[5])
);

DFFPOSX1 _1154_ (
    .CLK(clk_bF$buf5),
    .D(_40_),
    .Q(_589_[6])
);

DFFPOSX1 _1155_ (
    .CLK(clk_bF$buf4),
    .D(_41_),
    .Q(_589_[7])
);

DFFPOSX1 _1156_ (
    .CLK(clk_bF$buf3),
    .D(_42_),
    .Q(_589_[8])
);

DFFPOSX1 _1157_ (
    .CLK(clk_bF$buf2),
    .D(_43_),
    .Q(_589_[9])
);

DFFPOSX1 _1158_ (
    .CLK(clk_bF$buf1),
    .D(_44_),
    .Q(_589_[10])
);

DFFPOSX1 _1159_ (
    .CLK(clk_bF$buf0),
    .D(_45_),
    .Q(_589_[11])
);

DFFPOSX1 _1160_ (
    .CLK(clk_bF$buf8),
    .D(_46_),
    .Q(_589_[12])
);

DFFPOSX1 _1161_ (
    .CLK(clk_bF$buf7),
    .D(_47_),
    .Q(_589_[13])
);

DFFPOSX1 _1162_ (
    .CLK(clk_bF$buf6),
    .D(_48_),
    .Q(_589_[14])
);

DFFPOSX1 _1163_ (
    .CLK(clk_bF$buf5),
    .D(_49_),
    .Q(_589_[15])
);

DFFPOSX1 _1164_ (
    .CLK(clk_bF$buf4),
    .D(_50_),
    .Q(_589_[16])
);

DFFPOSX1 _1165_ (
    .CLK(clk_bF$buf3),
    .D(_51_),
    .Q(_589_[17])
);

DFFPOSX1 _1166_ (
    .CLK(clk_bF$buf2),
    .D(_52_),
    .Q(_589_[18])
);

DFFPOSX1 _1167_ (
    .CLK(clk_bF$buf1),
    .D(_53_),
    .Q(_589_[19])
);

DFFPOSX1 _1168_ (
    .CLK(clk_bF$buf0),
    .D(_54_),
    .Q(_589_[20])
);

DFFPOSX1 _1169_ (
    .CLK(clk_bF$buf8),
    .D(_55_),
    .Q(_589_[21])
);

DFFPOSX1 _1170_ (
    .CLK(clk_bF$buf7),
    .D(_56_),
    .Q(_589_[22])
);

DFFPOSX1 _1171_ (
    .CLK(clk_bF$buf6),
    .D(_57_),
    .Q(_589_[23])
);

DFFPOSX1 _1172_ (
    .CLK(clk_bF$buf5),
    .D(_58_),
    .Q(_590_[0])
);

DFFPOSX1 _1173_ (
    .CLK(clk_bF$buf4),
    .D(_59_),
    .Q(_590_[1])
);

DFFPOSX1 _1174_ (
    .CLK(clk_bF$buf3),
    .D(_60_),
    .Q(_590_[2])
);

DFFPOSX1 _1175_ (
    .CLK(clk_bF$buf2),
    .D(_61_),
    .Q(_590_[3])
);

DFFPOSX1 _1176_ (
    .CLK(clk_bF$buf1),
    .D(_62_),
    .Q(_590_[4])
);

DFFPOSX1 _1177_ (
    .CLK(clk_bF$buf0),
    .D(_63_),
    .Q(_590_[5])
);

DFFPOSX1 _1178_ (
    .CLK(clk_bF$buf8),
    .D(_64_),
    .Q(_590_[6])
);

DFFPOSX1 _1179_ (
    .CLK(clk_bF$buf7),
    .D(_65_),
    .Q(_590_[7])
);

DFFSR _1180_ (
    .CLK(clk_bF$buf6),
    .D(_66_),
    .Q(_592_[0]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1181_ (
    .CLK(clk_bF$buf5),
    .D(_67_),
    .Q(_592_[1]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1182_ (
    .CLK(clk_bF$buf4),
    .D(_68_),
    .Q(_592_[2]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1183_ (
    .CLK(clk_bF$buf3),
    .D(_69_),
    .Q(_592_[3]),
    .R(_0__bF$buf0),
    .S(vdd)
);

DFFSR _1184_ (
    .CLK(clk_bF$buf2),
    .D(_70_),
    .Q(_592_[4]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1185_ (
    .CLK(clk_bF$buf1),
    .D(_71_),
    .Q(_592_[5]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1186_ (
    .CLK(clk_bF$buf0),
    .D(_72_),
    .Q(_592_[6]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1187_ (
    .CLK(clk_bF$buf8),
    .D(_73_),
    .Q(_592_[7]),
    .R(_0__bF$buf0),
    .S(vdd)
);

DFFSR _1188_ (
    .CLK(clk_bF$buf7),
    .D(_74_),
    .Q(_592_[8]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1189_ (
    .CLK(clk_bF$buf6),
    .D(_75_),
    .Q(_592_[9]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1190_ (
    .CLK(clk_bF$buf5),
    .D(_76_),
    .Q(_592_[10]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1191_ (
    .CLK(clk_bF$buf4),
    .D(_77_),
    .Q(_592_[11]),
    .R(_0__bF$buf0),
    .S(vdd)
);

DFFSR _1192_ (
    .CLK(clk_bF$buf3),
    .D(_78_),
    .Q(_592_[12]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1193_ (
    .CLK(clk_bF$buf2),
    .D(_79_),
    .Q(_592_[13]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1194_ (
    .CLK(clk_bF$buf1),
    .D(_80_),
    .Q(_592_[14]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1195_ (
    .CLK(clk_bF$buf0),
    .D(_81_),
    .Q(_592_[15]),
    .R(_0__bF$buf0),
    .S(vdd)
);

DFFSR _1196_ (
    .CLK(clk_bF$buf8),
    .D(_82_),
    .Q(_592_[16]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1197_ (
    .CLK(clk_bF$buf7),
    .D(_83_),
    .Q(_592_[17]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1198_ (
    .CLK(clk_bF$buf6),
    .D(_84_),
    .Q(_592_[18]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1199_ (
    .CLK(clk_bF$buf5),
    .D(_85_),
    .Q(_592_[19]),
    .R(_0__bF$buf0),
    .S(vdd)
);

DFFSR _1200_ (
    .CLK(clk_bF$buf4),
    .D(_86_),
    .Q(_592_[20]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1201_ (
    .CLK(clk_bF$buf3),
    .D(_87_),
    .Q(_592_[21]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1202_ (
    .CLK(clk_bF$buf2),
    .D(_88_),
    .Q(_592_[22]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1203_ (
    .CLK(clk_bF$buf1),
    .D(_89_),
    .Q(_592_[23]),
    .R(_0__bF$buf0),
    .S(vdd)
);

INVX1 _1204_ (
    .A(\ALU_H4.a [0]),
    .Y(_525_)
);

INVX2 _1205_ (
    .A(instr[5]),
    .Y(_526_)
);

OAI21X1 _1206_ (
    .A(_526_),
    .B(\ALU_H4.b [0]),
    .C(_525_),
    .Y(_527_)
);

AOI21X1 _1207_ (
    .A(instr[4]),
    .B(\ALU_H4.b [0]),
    .C(_527_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_121 )
);

INVX1 _1208_ (
    .A(\ALU_H4.a [1]),
    .Y(_528_)
);

OAI21X1 _1209_ (
    .A(_526_),
    .B(\ALU_H4.b [1]),
    .C(_528_),
    .Y(_529_)
);

AOI21X1 _1210_ (
    .A(instr[4]),
    .B(\ALU_H4.b [1]),
    .C(_529_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_123 )
);

INVX1 _1211_ (
    .A(\ALU_H4.a [2]),
    .Y(_530_)
);

OAI21X1 _1212_ (
    .A(_526_),
    .B(\ALU_H4.b [2]),
    .C(_530_),
    .Y(_531_)
);

AOI21X1 _1213_ (
    .A(instr[4]),
    .B(\ALU_H4.b [2]),
    .C(_531_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_10 )
);

INVX2 _1214_ (
    .A(instr[7]),
    .Y(_532_)
);

AOI21X1 _1215_ (
    .A(\ALU_H4.b [0]),
    .B(_532_),
    .C(_525_),
    .Y(_533_)
);

OAI21X1 _1216_ (
    .A(\ALU_H4.b [0]),
    .B(instr[6]),
    .C(_533_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_120 )
);

AOI21X1 _1217_ (
    .A(\ALU_H4.b [1]),
    .B(_532_),
    .C(_528_),
    .Y(_534_)
);

OAI21X1 _1218_ (
    .A(\ALU_H4.b [1]),
    .B(instr[6]),
    .C(_534_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_122 )
);

AOI21X1 _1219_ (
    .A(\ALU_H4.b [2]),
    .B(_532_),
    .C(_530_),
    .Y(_535_)
);

OAI21X1 _1220_ (
    .A(\ALU_H4.b [2]),
    .B(instr[6]),
    .C(_535_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_11 )
);

INVX1 _1221_ (
    .A(\ALU_H4.a [3]),
    .Y(_536_)
);

OAI21X1 _1222_ (
    .A(_526_),
    .B(\ALU_H4.b [3]),
    .C(_536_),
    .Y(_537_)
);

AOI21X1 _1223_ (
    .A(instr[4]),
    .B(\ALU_H4.b [3]),
    .C(_537_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_127 )
);

AOI21X1 _1224_ (
    .A(\ALU_H4.b [3]),
    .B(_532_),
    .C(_536_),
    .Y(_538_)
);

OAI21X1 _1225_ (
    .A(instr[6]),
    .B(\ALU_H4.b [3]),
    .C(_538_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_126 )
);

NAND3X1 _1226_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_122 ),
    .B(\ALU_H4.SYNTHESIZED_WIRE_126 ),
    .C(\ALU_H4.SYNTHESIZED_WIRE_11 ),
    .Y(_539_)
);

INVX1 _1227_ (
    .A(_539_),
    .Y(_540_)
);

NAND2X1 _1228_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_120 ),
    .B(_540_),
    .Y(\ALU_H4.p )
);

INVX1 _1229_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_10 ),
    .Y(_541_)
);

NAND2X1 _1230_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_11 ),
    .B(\ALU_H4.SYNTHESIZED_WIRE_123 ),
    .Y(_542_)
);

NAND2X1 _1231_ (
    .A(_541_),
    .B(_542_),
    .Y(_543_)
);

INVX1 _1232_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_127 ),
    .Y(_544_)
);

INVX1 _1233_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_121 ),
    .Y(_545_)
);

OAI21X1 _1234_ (
    .A(_539_),
    .B(_545_),
    .C(_544_),
    .Y(_546_)
);

AOI21X1 _1235_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_126 ),
    .B(_543_),
    .C(_546_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_96 )
);

NOR2X1 _1236_ (
    .A(instr[3]),
    .B(_541_),
    .Y(_547_)
);

INVX2 _1237_ (
    .A(instr[3]),
    .Y(_548_)
);

NAND2X1 _1238_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_123 ),
    .B(_548_),
    .Y(_549_)
);

NAND3X1 _1239_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_122 ),
    .B(\ALU_H4.SYNTHESIZED_WIRE_121 ),
    .C(_548_),
    .Y(_550_)
);

AND2X2 _1240_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_120 ),
    .B(instr[2]),
    .Y(_551_)
);

NAND3X1 _1241_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_122 ),
    .B(_548_),
    .C(_551_),
    .Y(_552_)
);

NAND3X1 _1242_ (
    .A(_549_),
    .B(_550_),
    .C(_552_),
    .Y(_553_)
);

AOI21X1 _1243_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_11 ),
    .B(_553_),
    .C(_547_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_93 )
);

INVX1 _1244_ (
    .A(_553_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_106 )
);

INVX1 _1245_ (
    .A(instr[2]),
    .Y(_554_)
);

OAI21X1 _1246_ (
    .A(_554_),
    .B(\ALU_H4.p ),
    .C(\ALU_H4.SYNTHESIZED_WIRE_96 ),
    .Y(\ALU_H4.cout )
);

NOR2X1 _1247_ (
    .A(instr[3]),
    .B(_554_),
    .Y(_555_)
);

AOI22X1 _1248_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_121 ),
    .B(_548_),
    .C(_555_),
    .D(\ALU_H4.SYNTHESIZED_WIRE_120 ),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_104 )
);

XNOR2X1 _1249_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_126 ),
    .B(\ALU_H4.SYNTHESIZED_WIRE_93 ),
    .Y(_556_)
);

XNOR2X1 _1250_ (
    .A(_556_),
    .B(\ALU_H4.SYNTHESIZED_WIRE_127 ),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_107 )
);

XOR2X1 _1251_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_120 ),
    .B(\ALU_H4.SYNTHESIZED_WIRE_121 ),
    .Y(_557_)
);

XNOR2X1 _1252_ (
    .A(_557_),
    .B(_555_),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_110 )
);

XNOR2X1 _1253_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_122 ),
    .B(\ALU_H4.SYNTHESIZED_WIRE_104 ),
    .Y(_558_)
);

XNOR2X1 _1254_ (
    .A(_558_),
    .B(\ALU_H4.SYNTHESIZED_WIRE_123 ),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_109 )
);

XNOR2X1 _1255_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_11 ),
    .B(\ALU_H4.SYNTHESIZED_WIRE_106 ),
    .Y(_522_)
);

XNOR2X1 _1256_ (
    .A(_522_),
    .B(\ALU_H4.SYNTHESIZED_WIRE_10 ),
    .Y(\ALU_H4.SYNTHESIZED_WIRE_108 )
);

NAND2X1 _1257_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_108 ),
    .B(\ALU_H4.SYNTHESIZED_WIRE_107 ),
    .Y(_523_)
);

NAND2X1 _1258_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_109 ),
    .B(\ALU_H4.SYNTHESIZED_WIRE_110 ),
    .Y(_524_)
);

NOR2X1 _1259_ (
    .A(_523_),
    .B(_524_),
    .Y(\ALU_H4.eqv )
);

INVX1 _1260_ (
    .A(\ALU_L4.a [0]),
    .Y(_562_)
);

INVX2 _1261_ (
    .A(instr[5]),
    .Y(_563_)
);

OAI21X1 _1262_ (
    .A(_563_),
    .B(\ALU_L4.b [0]),
    .C(_562_),
    .Y(_564_)
);

AOI21X1 _1263_ (
    .A(instr[4]),
    .B(\ALU_L4.b [0]),
    .C(_564_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_121 )
);

INVX1 _1264_ (
    .A(\ALU_L4.a [1]),
    .Y(_565_)
);

OAI21X1 _1265_ (
    .A(_563_),
    .B(\ALU_L4.b [1]),
    .C(_565_),
    .Y(_566_)
);

AOI21X1 _1266_ (
    .A(instr[4]),
    .B(\ALU_L4.b [1]),
    .C(_566_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_123 )
);

INVX1 _1267_ (
    .A(\ALU_L4.a [2]),
    .Y(_567_)
);

OAI21X1 _1268_ (
    .A(_563_),
    .B(\ALU_L4.b [2]),
    .C(_567_),
    .Y(_568_)
);

AOI21X1 _1269_ (
    .A(instr[4]),
    .B(\ALU_L4.b [2]),
    .C(_568_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_10 )
);

INVX2 _1270_ (
    .A(instr[7]),
    .Y(_569_)
);

AOI21X1 _1271_ (
    .A(\ALU_L4.b [0]),
    .B(_569_),
    .C(_562_),
    .Y(_570_)
);

OAI21X1 _1272_ (
    .A(\ALU_L4.b [0]),
    .B(instr[6]),
    .C(_570_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_120 )
);

AOI21X1 _1273_ (
    .A(\ALU_L4.b [1]),
    .B(_569_),
    .C(_565_),
    .Y(_571_)
);

OAI21X1 _1274_ (
    .A(\ALU_L4.b [1]),
    .B(instr[6]),
    .C(_571_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_122 )
);

AOI21X1 _1275_ (
    .A(\ALU_L4.b [2]),
    .B(_569_),
    .C(_567_),
    .Y(_572_)
);

OAI21X1 _1276_ (
    .A(\ALU_L4.b [2]),
    .B(instr[6]),
    .C(_572_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_11 )
);

INVX1 _1277_ (
    .A(\ALU_L4.a [3]),
    .Y(_573_)
);

OAI21X1 _1278_ (
    .A(_563_),
    .B(\ALU_L4.b [3]),
    .C(_573_),
    .Y(_574_)
);

AOI21X1 _1279_ (
    .A(instr[4]),
    .B(\ALU_L4.b [3]),
    .C(_574_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_127 )
);

AOI21X1 _1280_ (
    .A(\ALU_L4.b [3]),
    .B(_569_),
    .C(_573_),
    .Y(_575_)
);

OAI21X1 _1281_ (
    .A(instr[6]),
    .B(\ALU_L4.b [3]),
    .C(_575_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_126 )
);

INVX1 _1282_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_10 ),
    .Y(_576_)
);

NOR2X1 _1283_ (
    .A(instr[3]),
    .B(_576_),
    .Y(_577_)
);

INVX2 _1284_ (
    .A(instr[3]),
    .Y(_578_)
);

NAND2X1 _1285_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_123 ),
    .B(_578_),
    .Y(_579_)
);

NAND3X1 _1286_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_122 ),
    .B(\ALU_L4.SYNTHESIZED_WIRE_121 ),
    .C(_578_),
    .Y(_580_)
);

AND2X2 _1287_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_120 ),
    .B(instr[2]),
    .Y(_581_)
);

NAND3X1 _1288_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_122 ),
    .B(_578_),
    .C(_581_),
    .Y(_582_)
);

NAND3X1 _1289_ (
    .A(_579_),
    .B(_580_),
    .C(_582_),
    .Y(_583_)
);

AOI21X1 _1290_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_11 ),
    .B(_583_),
    .C(_577_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_93 )
);

INVX1 _1291_ (
    .A(_583_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_106 )
);

INVX1 _1292_ (
    .A(instr[2]),
    .Y(_584_)
);

NOR2X1 _1293_ (
    .A(instr[3]),
    .B(_584_),
    .Y(_585_)
);

AOI22X1 _1294_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_121 ),
    .B(_578_),
    .C(_585_),
    .D(\ALU_L4.SYNTHESIZED_WIRE_120 ),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_104 )
);

XNOR2X1 _1295_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_126 ),
    .B(\ALU_L4.SYNTHESIZED_WIRE_93 ),
    .Y(_586_)
);

XNOR2X1 _1296_ (
    .A(_586_),
    .B(\ALU_L4.SYNTHESIZED_WIRE_127 ),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_107 )
);

XOR2X1 _1297_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_120 ),
    .B(\ALU_L4.SYNTHESIZED_WIRE_121 ),
    .Y(_587_)
);

XNOR2X1 _1298_ (
    .A(_587_),
    .B(_585_),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_110 )
);

XNOR2X1 _1299_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_122 ),
    .B(\ALU_L4.SYNTHESIZED_WIRE_104 ),
    .Y(_588_)
);

XNOR2X1 _1300_ (
    .A(_588_),
    .B(\ALU_L4.SYNTHESIZED_WIRE_123 ),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_109 )
);

XNOR2X1 _1301_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_11 ),
    .B(\ALU_L4.SYNTHESIZED_WIRE_106 ),
    .Y(_559_)
);

XNOR2X1 _1302_ (
    .A(_559_),
    .B(\ALU_L4.SYNTHESIZED_WIRE_10 ),
    .Y(\ALU_L4.SYNTHESIZED_WIRE_108 )
);

NAND2X1 _1303_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_108 ),
    .B(\ALU_L4.SYNTHESIZED_WIRE_107 ),
    .Y(_560_)
);

NAND2X1 _1304_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_109 ),
    .B(\ALU_L4.SYNTHESIZED_WIRE_110 ),
    .Y(_561_)
);

NOR2X1 _1305_ (
    .A(_560_),
    .B(_561_),
    .Y(\ALU_L4.eqv )
);

BUFX2 _1306_ (
    .A(_589_[0]),
    .Y(daddr[0])
);

BUFX2 _1307_ (
    .A(_589_[1]),
    .Y(daddr[1])
);

BUFX2 _1308_ (
    .A(_589_[10]),
    .Y(daddr[10])
);

BUFX2 _1309_ (
    .A(_589_[11]),
    .Y(daddr[11])
);

BUFX2 _1310_ (
    .A(_589_[12]),
    .Y(daddr[12])
);

BUFX2 _1311_ (
    .A(_589_[13]),
    .Y(daddr[13])
);

BUFX2 _1312_ (
    .A(_589_[14]),
    .Y(daddr[14])
);

BUFX2 _1313_ (
    .A(_589_[15]),
    .Y(daddr[15])
);

BUFX2 _1314_ (
    .A(_589_[16]),
    .Y(daddr[16])
);

BUFX2 _1315_ (
    .A(_589_[17]),
    .Y(daddr[17])
);

BUFX2 _1316_ (
    .A(_589_[18]),
    .Y(daddr[18])
);

BUFX2 _1317_ (
    .A(_589_[19]),
    .Y(daddr[19])
);

BUFX2 _1318_ (
    .A(_589_[2]),
    .Y(daddr[2])
);

BUFX2 _1319_ (
    .A(_589_[20]),
    .Y(daddr[20])
);

BUFX2 _1320_ (
    .A(_589_[21]),
    .Y(daddr[21])
);

BUFX2 _1321_ (
    .A(_589_[22]),
    .Y(daddr[22])
);

BUFX2 _1322_ (
    .A(_589_[23]),
    .Y(daddr[23])
);

BUFX2 _1323_ (
    .A(_589_[3]),
    .Y(daddr[3])
);

BUFX2 _1324_ (
    .A(_589_[4]),
    .Y(daddr[4])
);

BUFX2 _1325_ (
    .A(_589_[5]),
    .Y(daddr[5])
);

BUFX2 _1326_ (
    .A(_589_[6]),
    .Y(daddr[6])
);

BUFX2 _1327_ (
    .A(_589_[7]),
    .Y(daddr[7])
);

BUFX2 _1328_ (
    .A(_589_[8]),
    .Y(daddr[8])
);

BUFX2 _1329_ (
    .A(_589_[9]),
    .Y(daddr[9])
);

BUFX2 _1330_ (
    .A(_590_[0]),
    .Y(ddata_o[0])
);

BUFX2 _1331_ (
    .A(_590_[1]),
    .Y(ddata_o[1])
);

BUFX2 _1332_ (
    .A(_590_[2]),
    .Y(ddata_o[2])
);

BUFX2 _1333_ (
    .A(_590_[3]),
    .Y(ddata_o[3])
);

BUFX2 _1334_ (
    .A(_590_[4]),
    .Y(ddata_o[4])
);

BUFX2 _1335_ (
    .A(_590_[5]),
    .Y(ddata_o[5])
);

BUFX2 _1336_ (
    .A(_590_[6]),
    .Y(ddata_o[6])
);

BUFX2 _1337_ (
    .A(_590_[7]),
    .Y(ddata_o[7])
);

BUFX2 _1338_ (
    .A(_591_),
    .Y(dwrite)
);

BUFX2 _1339_ (
    .A(_592_[0]),
    .Y(iaddr[0])
);

BUFX2 _1340_ (
    .A(_592_[1]),
    .Y(iaddr[1])
);

BUFX2 _1341_ (
    .A(_592_[10]),
    .Y(iaddr[10])
);

BUFX2 _1342_ (
    .A(_592_[11]),
    .Y(iaddr[11])
);

BUFX2 _1343_ (
    .A(_592_[12]),
    .Y(iaddr[12])
);

BUFX2 _1344_ (
    .A(_592_[13]),
    .Y(iaddr[13])
);

BUFX2 _1345_ (
    .A(_592_[14]),
    .Y(iaddr[14])
);

BUFX2 _1346_ (
    .A(_592_[15]),
    .Y(iaddr[15])
);

BUFX2 _1347_ (
    .A(_592_[16]),
    .Y(iaddr[16])
);

BUFX2 _1348_ (
    .A(_592_[17]),
    .Y(iaddr[17])
);

BUFX2 _1349_ (
    .A(_592_[18]),
    .Y(iaddr[18])
);

BUFX2 _1350_ (
    .A(_592_[19]),
    .Y(iaddr[19])
);

BUFX2 _1351_ (
    .A(_592_[2]),
    .Y(iaddr[2])
);

BUFX2 _1352_ (
    .A(_592_[20]),
    .Y(iaddr[20])
);

BUFX2 _1353_ (
    .A(_592_[21]),
    .Y(iaddr[21])
);

BUFX2 _1354_ (
    .A(_592_[22]),
    .Y(iaddr[22])
);

BUFX2 _1355_ (
    .A(_592_[23]),
    .Y(iaddr[23])
);

BUFX2 _1356_ (
    .A(_592_[3]),
    .Y(iaddr[3])
);

BUFX2 _1357_ (
    .A(_592_[4]),
    .Y(iaddr[4])
);

BUFX2 _1358_ (
    .A(_592_[5]),
    .Y(iaddr[5])
);

BUFX2 _1359_ (
    .A(_592_[6]),
    .Y(iaddr[6])
);

BUFX2 _1360_ (
    .A(_592_[7]),
    .Y(iaddr[7])
);

BUFX2 _1361_ (
    .A(_592_[8]),
    .Y(iaddr[8])
);

BUFX2 _1362_ (
    .A(_592_[9]),
    .Y(iaddr[9])
);

INVX8 _593_ (
    .A(rst),
    .Y(_0_)
);

INVX1 _594_ (
    .A(instr[13]),
    .Y(_90_)
);

INVX2 _595_ (
    .A(instr[14]),
    .Y(_91_)
);

AOI21X1 _596_ (
    .A(_90_),
    .B(_91_),
    .C(WAIT_bF$buf1),
    .Y(_92_)
);

INVX8 _597_ (
    .A(WAIT_bF$buf0),
    .Y(_93_)
);

NAND3X1 _598_ (
    .A(instr[13]),
    .B(instr[14]),
    .C(_93__bF$buf2),
    .Y(_94_)
);

INVX2 _599_ (
    .A(instr[15]),
    .Y(_95_)
);

NOR2X1 _600_ (
    .A(WAIT_bF$buf4),
    .B(instr[12]),
    .Y(_96_)
);

NAND3X1 _601_ (
    .A(instr[11]),
    .B(_95_),
    .C(_96_),
    .Y(_97_)
);

NOR2X1 _602_ (
    .A(instr[11]),
    .B(instr[12]),
    .Y(_98_)
);

NAND3X1 _603_ (
    .A(_93__bF$buf1),
    .B(instr[15]),
    .C(_98_),
    .Y(_99_)
);

OAI22X1 _604_ (
    .A(_97_),
    .B(_94_),
    .C(_92_),
    .D(_99_),
    .Y(_100_)
);

NAND3X1 _605_ (
    .A(instr[13]),
    .B(_93__bF$buf0),
    .C(_91_),
    .Y(_101_)
);

OAI21X1 _606_ (
    .A(instr[13]),
    .B(instr[14]),
    .C(_93__bF$buf4),
    .Y(_102_)
);

INVX1 _607_ (
    .A(instr[12]),
    .Y(_103_)
);

NOR3X1 _608_ (
    .A(instr[11]),
    .B(WAIT_bF$buf3),
    .C(_103_),
    .Y(_104_)
);

NAND3X1 _609_ (
    .A(instr[15]),
    .B(_102_),
    .C(_104_),
    .Y(_105_)
);

OAI21X1 _610_ (
    .A(_101_),
    .B(_99_),
    .C(_105_),
    .Y(_106_)
);

NOR2X1 _611_ (
    .A(_100_),
    .B(_106_),
    .Y(_107_)
);

NOR3X1 _612_ (
    .A(WAIT_bF$buf2),
    .B(instr[13]),
    .C(_91_),
    .Y(_108_)
);

NAND3X1 _613_ (
    .A(instr[15]),
    .B(_104_),
    .C(_108_),
    .Y(_109_)
);

OR2X2 _614_ (
    .A(_99_),
    .B(_94_),
    .Y(_110_)
);

AND2X2 _615_ (
    .A(_110_),
    .B(_109_),
    .Y(_111_)
);

NOR2X1 _616_ (
    .A(WAIT_bF$buf1),
    .B(_95_),
    .Y(_112_)
);

NAND2X1 _617_ (
    .A(instr[15]),
    .B(_93__bF$buf3),
    .Y(_113_)
);

INVX1 _618_ (
    .A(instr[11]),
    .Y(_114_)
);

NAND3X1 _619_ (
    .A(instr[12]),
    .B(_114_),
    .C(_93__bF$buf2),
    .Y(_115_)
);

NOR3X1 _620_ (
    .A(_115_),
    .B(_113_),
    .C(_101_),
    .Y(_116_)
);

OAI21X1 _621_ (
    .A(instr[11]),
    .B(instr[12]),
    .C(_93__bF$buf1),
    .Y(_117_)
);

AND2X2 _622_ (
    .A(_108_),
    .B(_117_),
    .Y(_118_)
);

AOI21X1 _623_ (
    .A(_112_),
    .B(_118_),
    .C(_116_),
    .Y(_119_)
);

NAND3X1 _624_ (
    .A(_111_),
    .B(_119_),
    .C(_107_),
    .Y(_120_)
);

NOR3X1 _625_ (
    .A(_115_),
    .B(_112_),
    .C(_92_),
    .Y(_121_)
);

INVX1 _626_ (
    .A(_121_),
    .Y(_122_)
);

OAI21X1 _627_ (
    .A(instr[15]),
    .B(_101_),
    .C(_122_),
    .Y(_123_)
);

INVX2 _628_ (
    .A(instr[9]),
    .Y(_124_)
);

NAND2X1 _629_ (
    .A(instr[8]),
    .B(_124_),
    .Y(_125_)
);

NOR2X1 _630_ (
    .A(instr[10]),
    .B(_125_),
    .Y(_126_)
);

OAI21X1 _631_ (
    .A(_120_),
    .B(_123_),
    .C(_126_),
    .Y(_127_)
);

NOR3X1 _632_ (
    .A(WAIT_bF$buf0),
    .B(instr[14]),
    .C(_90_),
    .Y(_128_)
);

NAND3X1 _633_ (
    .A(_112_),
    .B(_104_),
    .C(_128_),
    .Y(_129_)
);

NAND3X1 _634_ (
    .A(_112_),
    .B(_117_),
    .C(_128_),
    .Y(_130_)
);

AND2X2 _635_ (
    .A(_105_),
    .B(_130_),
    .Y(_131_)
);

NAND3X1 _636_ (
    .A(instr[11]),
    .B(instr[12]),
    .C(_93__bF$buf0),
    .Y(_132_)
);

NOR3X1 _637_ (
    .A(_132_),
    .B(_112_),
    .C(_101_),
    .Y(_133_)
);

NOR2X1 _638_ (
    .A(_133_),
    .B(_100_),
    .Y(_134_)
);

NAND3X1 _639_ (
    .A(_129_),
    .B(_131_),
    .C(_134_),
    .Y(_135_)
);

NAND3X1 _640_ (
    .A(instr[14]),
    .B(_117_),
    .C(_112_),
    .Y(_136_)
);

AND2X2 _641_ (
    .A(_109_),
    .B(_136_),
    .Y(_137_)
);

NAND3X1 _642_ (
    .A(_95_),
    .B(_104_),
    .C(_128_),
    .Y(_138_)
);

NAND3X1 _643_ (
    .A(_95_),
    .B(_117_),
    .C(_128_),
    .Y(_139_)
);

AND2X2 _644_ (
    .A(_138_),
    .B(_139_),
    .Y(_140_)
);

NAND3X1 _645_ (
    .A(_122_),
    .B(_137_),
    .C(_140_),
    .Y(_141_)
);

NOR2X1 _646_ (
    .A(_141_),
    .B(_135_),
    .Y(_142_)
);

OAI21X1 _647_ (
    .A(_91_),
    .B(_99_),
    .C(_109_),
    .Y(_143_)
);

NAND2X1 _648_ (
    .A(\ALU_L4.b [1]),
    .B(_143_),
    .Y(_144_)
);

AOI22X1 _649_ (
    .A(\ALU_L4.SYNTHESIZED_WIRE_110 ),
    .B(_121_),
    .C(_106_),
    .D(\ALU_L4.a [1]),
    .Y(_145_)
);

INVX1 _650_ (
    .A(D[0]),
    .Y(_146_)
);

INVX1 _651_ (
    .A(ddata_i[0]),
    .Y(_147_)
);

NOR2X1 _652_ (
    .A(WAIT_bF$buf4),
    .B(_103_),
    .Y(_148_)
);

NOR2X1 _653_ (
    .A(instr[15]),
    .B(_114_),
    .Y(_149_)
);

NAND3X1 _654_ (
    .A(_148_),
    .B(_149_),
    .C(_128_),
    .Y(_150_)
);

OAI22X1 _655_ (
    .A(_150_),
    .B(_146_),
    .C(_147_),
    .D(_139_),
    .Y(_151_)
);

INVX2 _656_ (
    .A(\ALU_H4.b [3]),
    .Y(_152_)
);

INVX1 _657_ (
    .A(instr[0]),
    .Y(_153_)
);

NAND3X1 _658_ (
    .A(_102_),
    .B(_117_),
    .C(_112_),
    .Y(_154_)
);

OAI22X1 _659_ (
    .A(_152_),
    .B(_154_),
    .C(_138_),
    .D(_153_),
    .Y(_155_)
);

NOR2X1 _660_ (
    .A(_151_),
    .B(_155_),
    .Y(_156_)
);

NAND3X1 _661_ (
    .A(_144_),
    .B(_145_),
    .C(_156_),
    .Y(_157_)
);

AOI21X1 _662_ (
    .A(C[0]),
    .B(_142_),
    .C(_157_),
    .Y(_158_)
);

OR2X2 _663_ (
    .A(_106_),
    .B(_100_),
    .Y(_159_)
);

NAND2X1 _664_ (
    .A(_119_),
    .B(_111_),
    .Y(_160_)
);

NOR3X1 _665_ (
    .A(_159_),
    .B(_123_),
    .C(_160_),
    .Y(_161_)
);

INVX4 _666_ (
    .A(_126_),
    .Y(_162_)
);

OAI21X1 _667_ (
    .A(_161__bF$buf7),
    .B(_162_),
    .C(\ALU_L4.a [0]),
    .Y(_163_)
);

OAI21X1 _668_ (
    .A(_158_),
    .B(_127_),
    .C(_163_),
    .Y(_1_)
);

AOI22X1 _669_ (
    .A(\ALU_L4.b [0]),
    .B(_116_),
    .C(_100_),
    .D(\ALU_L4.a [0]),
    .Y(_164_)
);

AOI22X1 _670_ (
    .A(_133_),
    .B(D[1]),
    .C(\ALU_L4.SYNTHESIZED_WIRE_109 ),
    .D(_121_),
    .Y(_165_)
);

AND2X2 _671_ (
    .A(_164_),
    .B(_165_),
    .Y(_166_)
);

INVX1 _672_ (
    .A(\ALU_L4.a [2]),
    .Y(_167_)
);

AOI21X1 _673_ (
    .A(_105_),
    .B(_130_),
    .C(_167_),
    .Y(_168_)
);

INVX1 _674_ (
    .A(\ALU_L4.b [2]),
    .Y(_169_)
);

AOI21X1 _675_ (
    .A(_136_),
    .B(_109_),
    .C(_169_),
    .Y(_170_)
);

INVX1 _676_ (
    .A(instr[1]),
    .Y(_171_)
);

INVX1 _677_ (
    .A(ddata_i[1]),
    .Y(_172_)
);

OAI22X1 _678_ (
    .A(_139_),
    .B(_172_),
    .C(_138_),
    .D(_171_),
    .Y(_173_)
);

NOR3X1 _679_ (
    .A(_170_),
    .B(_168_),
    .C(_173_),
    .Y(_174_)
);

NAND2X1 _680_ (
    .A(_166_),
    .B(_174_),
    .Y(_175_)
);

AOI21X1 _681_ (
    .A(C[1]),
    .B(_142_),
    .C(_175_),
    .Y(_176_)
);

OAI21X1 _682_ (
    .A(_161__bF$buf6),
    .B(_162_),
    .C(\ALU_L4.a [1]),
    .Y(_177_)
);

OAI21X1 _683_ (
    .A(_176_),
    .B(_127_),
    .C(_177_),
    .Y(_2_)
);

AOI22X1 _684_ (
    .A(_121_),
    .B(\ALU_L4.SYNTHESIZED_WIRE_108 ),
    .C(\ALU_L4.b [1]),
    .D(_116_),
    .Y(_178_)
);

AOI22X1 _685_ (
    .A(D[2]),
    .B(_133_),
    .C(_100_),
    .D(\ALU_L4.a [1]),
    .Y(_179_)
);

AND2X2 _686_ (
    .A(_179_),
    .B(_178_),
    .Y(_180_)
);

INVX1 _687_ (
    .A(\ALU_L4.a [3]),
    .Y(_181_)
);

AOI21X1 _688_ (
    .A(_105_),
    .B(_130_),
    .C(_181_),
    .Y(_182_)
);

INVX1 _689_ (
    .A(\ALU_L4.b [3]),
    .Y(_183_)
);

AOI21X1 _690_ (
    .A(_136_),
    .B(_109_),
    .C(_183_),
    .Y(_184_)
);

INVX1 _691_ (
    .A(instr[2]),
    .Y(_185_)
);

INVX1 _692_ (
    .A(ddata_i[2]),
    .Y(_186_)
);

OAI22X1 _693_ (
    .A(_139_),
    .B(_186_),
    .C(_138_),
    .D(_185_),
    .Y(_187_)
);

NOR3X1 _694_ (
    .A(_184_),
    .B(_182_),
    .C(_187_),
    .Y(_188_)
);

NAND2X1 _695_ (
    .A(_188_),
    .B(_180_),
    .Y(_189_)
);

AOI21X1 _696_ (
    .A(C[2]),
    .B(_142_),
    .C(_189_),
    .Y(_190_)
);

OAI21X1 _697_ (
    .A(_161__bF$buf5),
    .B(_162_),
    .C(\ALU_L4.a [2]),
    .Y(_191_)
);

OAI21X1 _698_ (
    .A(_190_),
    .B(_127_),
    .C(_191_),
    .Y(_3_)
);

AOI22X1 _699_ (
    .A(\ALU_L4.b [2]),
    .B(_116_),
    .C(_100_),
    .D(\ALU_L4.a [2]),
    .Y(_192_)
);

AOI22X1 _700_ (
    .A(_133_),
    .B(D[3]),
    .C(\ALU_L4.SYNTHESIZED_WIRE_107 ),
    .D(_121_),
    .Y(_193_)
);

AND2X2 _701_ (
    .A(_192_),
    .B(_193_),
    .Y(_194_)
);

INVX1 _702_ (
    .A(\ALU_H4.a [0]),
    .Y(_195_)
);

AOI21X1 _703_ (
    .A(_105_),
    .B(_130_),
    .C(_195_),
    .Y(_196_)
);

INVX1 _704_ (
    .A(\ALU_H4.b [0]),
    .Y(_197_)
);

AOI21X1 _705_ (
    .A(_136_),
    .B(_109_),
    .C(_197_),
    .Y(_198_)
);

INVX1 _706_ (
    .A(instr[3]),
    .Y(_199_)
);

INVX1 _707_ (
    .A(ddata_i[3]),
    .Y(_200_)
);

OAI22X1 _708_ (
    .A(_139_),
    .B(_200_),
    .C(_138_),
    .D(_199_),
    .Y(_201_)
);

NOR3X1 _709_ (
    .A(_198_),
    .B(_196_),
    .C(_201_),
    .Y(_202_)
);

NAND2X1 _710_ (
    .A(_194_),
    .B(_202_),
    .Y(_203_)
);

AOI21X1 _711_ (
    .A(C[3]),
    .B(_142_),
    .C(_203_),
    .Y(_204_)
);

OAI21X1 _712_ (
    .A(_161__bF$buf4),
    .B(_162_),
    .C(\ALU_L4.a [3]),
    .Y(_205_)
);

OAI21X1 _713_ (
    .A(_204_),
    .B(_127_),
    .C(_205_),
    .Y(_4_)
);

AOI22X1 _714_ (
    .A(\ALU_L4.b [3]),
    .B(_116_),
    .C(_100_),
    .D(\ALU_L4.a [3]),
    .Y(_206_)
);

AOI22X1 _715_ (
    .A(_133_),
    .B(D[4]),
    .C(\ALU_H4.SYNTHESIZED_WIRE_110 ),
    .D(_121_),
    .Y(_207_)
);

AND2X2 _716_ (
    .A(_206_),
    .B(_207_),
    .Y(_208_)
);

INVX1 _717_ (
    .A(\ALU_H4.a [1]),
    .Y(_209_)
);

AOI21X1 _718_ (
    .A(_105_),
    .B(_130_),
    .C(_209_),
    .Y(_210_)
);

INVX1 _719_ (
    .A(\ALU_H4.b [1]),
    .Y(_211_)
);

AOI21X1 _720_ (
    .A(_136_),
    .B(_109_),
    .C(_211_),
    .Y(_212_)
);

INVX1 _721_ (
    .A(instr[4]),
    .Y(_213_)
);

INVX1 _722_ (
    .A(ddata_i[4]),
    .Y(_214_)
);

OAI22X1 _723_ (
    .A(_139_),
    .B(_214_),
    .C(_138_),
    .D(_213_),
    .Y(_215_)
);

NOR3X1 _724_ (
    .A(_212_),
    .B(_210_),
    .C(_215_),
    .Y(_216_)
);

NAND2X1 _725_ (
    .A(_208_),
    .B(_216_),
    .Y(_217_)
);

AOI21X1 _726_ (
    .A(C[4]),
    .B(_142_),
    .C(_217_),
    .Y(_218_)
);

OAI21X1 _727_ (
    .A(_161__bF$buf3),
    .B(_162_),
    .C(\ALU_H4.a [0]),
    .Y(_219_)
);

OAI21X1 _728_ (
    .A(_218_),
    .B(_127_),
    .C(_219_),
    .Y(_5_)
);

AOI22X1 _729_ (
    .A(\ALU_H4.b [0]),
    .B(_116_),
    .C(_100_),
    .D(\ALU_H4.a [0]),
    .Y(_220_)
);

AOI22X1 _730_ (
    .A(_133_),
    .B(D[5]),
    .C(\ALU_H4.SYNTHESIZED_WIRE_109 ),
    .D(_121_),
    .Y(_221_)
);

AND2X2 _731_ (
    .A(_220_),
    .B(_221_),
    .Y(_222_)
);

INVX1 _732_ (
    .A(\ALU_H4.a [2]),
    .Y(_223_)
);

AOI21X1 _733_ (
    .A(_105_),
    .B(_130_),
    .C(_223_),
    .Y(_224_)
);

INVX1 _734_ (
    .A(\ALU_H4.b [2]),
    .Y(_225_)
);

AOI21X1 _735_ (
    .A(_136_),
    .B(_109_),
    .C(_225_),
    .Y(_226_)
);

INVX1 _736_ (
    .A(instr[5]),
    .Y(_227_)
);

INVX1 _737_ (
    .A(ddata_i[5]),
    .Y(_228_)
);

OAI22X1 _738_ (
    .A(_139_),
    .B(_228_),
    .C(_138_),
    .D(_227_),
    .Y(_229_)
);

NOR3X1 _739_ (
    .A(_226_),
    .B(_224_),
    .C(_229_),
    .Y(_230_)
);

NAND2X1 _740_ (
    .A(_222_),
    .B(_230_),
    .Y(_231_)
);

AOI21X1 _741_ (
    .A(C[5]),
    .B(_142_),
    .C(_231_),
    .Y(_232_)
);

OAI21X1 _742_ (
    .A(_161__bF$buf2),
    .B(_162_),
    .C(\ALU_H4.a [1]),
    .Y(_233_)
);

OAI21X1 _743_ (
    .A(_232_),
    .B(_127_),
    .C(_233_),
    .Y(_6_)
);

AOI22X1 _744_ (
    .A(\ALU_H4.b [1]),
    .B(_116_),
    .C(_100_),
    .D(\ALU_H4.a [1]),
    .Y(_234_)
);

AOI22X1 _745_ (
    .A(_133_),
    .B(D[6]),
    .C(\ALU_H4.SYNTHESIZED_WIRE_108 ),
    .D(_121_),
    .Y(_235_)
);

AND2X2 _746_ (
    .A(_234_),
    .B(_235_),
    .Y(_236_)
);

INVX2 _747_ (
    .A(\ALU_H4.a [3]),
    .Y(_237_)
);

AOI21X1 _748_ (
    .A(_105_),
    .B(_130_),
    .C(_237_),
    .Y(_238_)
);

AOI21X1 _749_ (
    .A(_136_),
    .B(_109_),
    .C(_152_),
    .Y(_239_)
);

INVX1 _750_ (
    .A(instr[6]),
    .Y(_240_)
);

INVX1 _751_ (
    .A(ddata_i[6]),
    .Y(_241_)
);

OAI22X1 _752_ (
    .A(_139_),
    .B(_241_),
    .C(_138_),
    .D(_240_),
    .Y(_242_)
);

NOR3X1 _753_ (
    .A(_239_),
    .B(_238_),
    .C(_242_),
    .Y(_243_)
);

NAND2X1 _754_ (
    .A(_236_),
    .B(_243_),
    .Y(_244_)
);

AOI21X1 _755_ (
    .A(C[6]),
    .B(_142_),
    .C(_244_),
    .Y(_245_)
);

OAI21X1 _756_ (
    .A(_161__bF$buf1),
    .B(_162_),
    .C(\ALU_H4.a [2]),
    .Y(_246_)
);

OAI21X1 _757_ (
    .A(_245_),
    .B(_127_),
    .C(_246_),
    .Y(_7_)
);

INVX1 _758_ (
    .A(instr[7]),
    .Y(_247_)
);

OAI22X1 _759_ (
    .A(_138_),
    .B(_247_),
    .C(_225_),
    .D(_129_),
    .Y(_248_)
);

INVX1 _760_ (
    .A(ddata_i[7]),
    .Y(_249_)
);

OAI22X1 _761_ (
    .A(_139_),
    .B(_249_),
    .C(_109_),
    .D(_152_),
    .Y(_250_)
);

NOR2X1 _762_ (
    .A(_250_),
    .B(_248_),
    .Y(_251_)
);

NAND3X1 _763_ (
    .A(\ALU_L4.a [0]),
    .B(_117_),
    .C(_112_),
    .Y(_252_)
);

OAI22X1 _764_ (
    .A(_94_),
    .B(_252_),
    .C(_130_),
    .D(_237_),
    .Y(_253_)
);

AOI21X1 _765_ (
    .A(D[7]),
    .B(_133_),
    .C(_253_),
    .Y(_254_)
);

AOI22X1 _766_ (
    .A(\ALU_H4.SYNTHESIZED_WIRE_107 ),
    .B(_121_),
    .C(_100_),
    .D(\ALU_H4.a [2]),
    .Y(_255_)
);

NAND3X1 _767_ (
    .A(_255_),
    .B(_254_),
    .C(_251_),
    .Y(_256_)
);

AOI21X1 _768_ (
    .A(C[7]),
    .B(_142_),
    .C(_256_),
    .Y(_257_)
);

OAI21X1 _769_ (
    .A(_161__bF$buf0),
    .B(_162_),
    .C(\ALU_H4.a [3]),
    .Y(_258_)
);

OAI21X1 _770_ (
    .A(_257_),
    .B(_127_),
    .C(_258_),
    .Y(_8_)
);

NOR3X1 _771_ (
    .A(instr[10]),
    .B(instr[8]),
    .C(_124_),
    .Y(_259_)
);

OAI21X1 _772_ (
    .A(_120_),
    .B(_123_),
    .C(_259_),
    .Y(_260_)
);

INVX4 _773_ (
    .A(_259_),
    .Y(_261_)
);

OAI21X1 _774_ (
    .A(_161__bF$buf7),
    .B(_261_),
    .C(\ALU_L4.b [0]),
    .Y(_262_)
);

OAI21X1 _775_ (
    .A(_158_),
    .B(_260_),
    .C(_262_),
    .Y(_9_)
);

OAI21X1 _776_ (
    .A(_161__bF$buf6),
    .B(_261_),
    .C(\ALU_L4.b [1]),
    .Y(_263_)
);

OAI21X1 _777_ (
    .A(_176_),
    .B(_260_),
    .C(_263_),
    .Y(_10_)
);

OAI21X1 _778_ (
    .A(_161__bF$buf5),
    .B(_261_),
    .C(\ALU_L4.b [2]),
    .Y(_264_)
);

OAI21X1 _779_ (
    .A(_190_),
    .B(_260_),
    .C(_264_),
    .Y(_11_)
);

OAI21X1 _780_ (
    .A(_161__bF$buf4),
    .B(_261_),
    .C(\ALU_L4.b [3]),
    .Y(_265_)
);

OAI21X1 _781_ (
    .A(_204_),
    .B(_260_),
    .C(_265_),
    .Y(_12_)
);

OAI21X1 _782_ (
    .A(_161__bF$buf3),
    .B(_261_),
    .C(\ALU_H4.b [0]),
    .Y(_266_)
);

OAI21X1 _783_ (
    .A(_218_),
    .B(_260_),
    .C(_266_),
    .Y(_13_)
);

OAI21X1 _784_ (
    .A(_161__bF$buf2),
    .B(_261_),
    .C(\ALU_H4.b [1]),
    .Y(_267_)
);

OAI21X1 _785_ (
    .A(_232_),
    .B(_260_),
    .C(_267_),
    .Y(_14_)
);

OAI21X1 _786_ (
    .A(_161__bF$buf1),
    .B(_261_),
    .C(\ALU_H4.b [2]),
    .Y(_268_)
);

OAI21X1 _787_ (
    .A(_245_),
    .B(_260_),
    .C(_268_),
    .Y(_15_)
);

OAI21X1 _788_ (
    .A(_161__bF$buf0),
    .B(_261_),
    .C(\ALU_H4.b [3]),
    .Y(_269_)
);

OAI21X1 _789_ (
    .A(_257_),
    .B(_260_),
    .C(_269_),
    .Y(_16_)
);

NOR2X1 _790_ (
    .A(instr[9]),
    .B(instr[8]),
    .Y(_270_)
);

INVX1 _791_ (
    .A(_270_),
    .Y(_271_)
);

NOR2X1 _792_ (
    .A(instr[10]),
    .B(_271_),
    .Y(_272_)
);

OAI21X1 _793_ (
    .A(_120_),
    .B(_123_),
    .C(_272_),
    .Y(_273_)
);

INVX4 _794_ (
    .A(_272_),
    .Y(_274_)
);

OAI21X1 _795_ (
    .A(_161__bF$buf7),
    .B(_274_),
    .C(C[0]),
    .Y(_275_)
);

OAI21X1 _796_ (
    .A(_158_),
    .B(_273_),
    .C(_275_),
    .Y(_17_)
);

OAI21X1 _797_ (
    .A(_161__bF$buf6),
    .B(_274_),
    .C(C[1]),
    .Y(_276_)
);

OAI21X1 _798_ (
    .A(_176_),
    .B(_273_),
    .C(_276_),
    .Y(_18_)
);

OAI21X1 _799_ (
    .A(_161__bF$buf5),
    .B(_274_),
    .C(C[2]),
    .Y(_277_)
);

OAI21X1 _800_ (
    .A(_190_),
    .B(_273_),
    .C(_277_),
    .Y(_19_)
);

OAI21X1 _801_ (
    .A(_161__bF$buf4),
    .B(_274_),
    .C(C[3]),
    .Y(_278_)
);

OAI21X1 _802_ (
    .A(_204_),
    .B(_273_),
    .C(_278_),
    .Y(_20_)
);

OAI21X1 _803_ (
    .A(_161__bF$buf3),
    .B(_274_),
    .C(C[4]),
    .Y(_279_)
);

OAI21X1 _804_ (
    .A(_218_),
    .B(_273_),
    .C(_279_),
    .Y(_21_)
);

OAI21X1 _805_ (
    .A(_161__bF$buf2),
    .B(_274_),
    .C(C[5]),
    .Y(_280_)
);

OAI21X1 _806_ (
    .A(_232_),
    .B(_273_),
    .C(_280_),
    .Y(_22_)
);

OAI21X1 _807_ (
    .A(_161__bF$buf1),
    .B(_274_),
    .C(C[6]),
    .Y(_281_)
);

OAI21X1 _808_ (
    .A(_245_),
    .B(_273_),
    .C(_281_),
    .Y(_23_)
);

OAI21X1 _809_ (
    .A(_161__bF$buf0),
    .B(_274_),
    .C(C[7]),
    .Y(_282_)
);

OAI21X1 _810_ (
    .A(_257_),
    .B(_273_),
    .C(_282_),
    .Y(_24_)
);

NOR2X1 _811_ (
    .A(instr[8]),
    .B(_124_),
    .Y(_283_)
);

NAND2X1 _812_ (
    .A(instr[10]),
    .B(_283_),
    .Y(_284_)
);

INVX1 _813_ (
    .A(_284_),
    .Y(_285_)
);

OAI21X1 _814_ (
    .A(_120_),
    .B(_123_),
    .C(_285_),
    .Y(_286_)
);

OAI21X1 _815_ (
    .A(_161__bF$buf7),
    .B(_284_),
    .C(D[0]),
    .Y(_287_)
);

OAI21X1 _816_ (
    .A(_158_),
    .B(_286_),
    .C(_287_),
    .Y(_25_)
);

OAI21X1 _817_ (
    .A(_161__bF$buf6),
    .B(_284_),
    .C(D[1]),
    .Y(_288_)
);

OAI21X1 _818_ (
    .A(_176_),
    .B(_286_),
    .C(_288_),
    .Y(_26_)
);

OAI21X1 _819_ (
    .A(_161__bF$buf5),
    .B(_284_),
    .C(D[2]),
    .Y(_289_)
);

OAI21X1 _820_ (
    .A(_190_),
    .B(_286_),
    .C(_289_),
    .Y(_27_)
);

OAI21X1 _821_ (
    .A(_161__bF$buf4),
    .B(_284_),
    .C(D[3]),
    .Y(_290_)
);

OAI21X1 _822_ (
    .A(_204_),
    .B(_286_),
    .C(_290_),
    .Y(_28_)
);

OAI21X1 _823_ (
    .A(_161__bF$buf3),
    .B(_284_),
    .C(D[4]),
    .Y(_291_)
);

OAI21X1 _824_ (
    .A(_218_),
    .B(_286_),
    .C(_291_),
    .Y(_29_)
);

OAI21X1 _825_ (
    .A(_161__bF$buf2),
    .B(_284_),
    .C(D[5]),
    .Y(_292_)
);

OAI21X1 _826_ (
    .A(_232_),
    .B(_286_),
    .C(_292_),
    .Y(_30_)
);

OAI21X1 _827_ (
    .A(_161__bF$buf1),
    .B(_284_),
    .C(D[6]),
    .Y(_293_)
);

OAI21X1 _828_ (
    .A(_245_),
    .B(_286_),
    .C(_293_),
    .Y(_31_)
);

OAI21X1 _829_ (
    .A(_161__bF$buf0),
    .B(_284_),
    .C(D[7]),
    .Y(_294_)
);

OAI21X1 _830_ (
    .A(_257_),
    .B(_286_),
    .C(_294_),
    .Y(_32_)
);

NAND2X1 _831_ (
    .A(instr[9]),
    .B(instr[8]),
    .Y(_295_)
);

NOR2X1 _832_ (
    .A(instr[10]),
    .B(_295_),
    .Y(_296_)
);

OAI21X1 _833_ (
    .A(_120_),
    .B(_123_),
    .C(_296_),
    .Y(_297_)
);

INVX4 _834_ (
    .A(_296_),
    .Y(_298_)
);

OAI21X1 _835_ (
    .A(_161__bF$buf7),
    .B(_298_),
    .C(_589_[0]),
    .Y(_299_)
);

OAI21X1 _836_ (
    .A(_158_),
    .B(_297_),
    .C(_299_),
    .Y(_34_)
);

OAI21X1 _837_ (
    .A(_161__bF$buf6),
    .B(_298_),
    .C(_589_[1]),
    .Y(_300_)
);

OAI21X1 _838_ (
    .A(_176_),
    .B(_297_),
    .C(_300_),
    .Y(_35_)
);

OAI21X1 _839_ (
    .A(_161__bF$buf5),
    .B(_298_),
    .C(_589_[2]),
    .Y(_301_)
);

OAI21X1 _840_ (
    .A(_190_),
    .B(_297_),
    .C(_301_),
    .Y(_36_)
);

OAI21X1 _841_ (
    .A(_161__bF$buf4),
    .B(_298_),
    .C(_589_[3]),
    .Y(_302_)
);

OAI21X1 _842_ (
    .A(_204_),
    .B(_297_),
    .C(_302_),
    .Y(_37_)
);

OAI21X1 _843_ (
    .A(_161__bF$buf3),
    .B(_298_),
    .C(_589_[4]),
    .Y(_303_)
);

OAI21X1 _844_ (
    .A(_218_),
    .B(_297_),
    .C(_303_),
    .Y(_38_)
);

OAI21X1 _845_ (
    .A(_161__bF$buf2),
    .B(_298_),
    .C(_589_[5]),
    .Y(_304_)
);

OAI21X1 _846_ (
    .A(_232_),
    .B(_297_),
    .C(_304_),
    .Y(_39_)
);

OAI21X1 _847_ (
    .A(_161__bF$buf1),
    .B(_298_),
    .C(_589_[6]),
    .Y(_305_)
);

OAI21X1 _848_ (
    .A(_245_),
    .B(_297_),
    .C(_305_),
    .Y(_40_)
);

OAI21X1 _849_ (
    .A(_161__bF$buf0),
    .B(_298_),
    .C(_589_[7]),
    .Y(_306_)
);

OAI21X1 _850_ (
    .A(_257_),
    .B(_297_),
    .C(_306_),
    .Y(_41_)
);

INVX2 _851_ (
    .A(instr[10]),
    .Y(_307_)
);

NOR2X1 _852_ (
    .A(_307_),
    .B(_271_),
    .Y(_308_)
);

OAI21X1 _853_ (
    .A(_120_),
    .B(_123_),
    .C(_308_),
    .Y(_309_)
);

INVX4 _854_ (
    .A(_308_),
    .Y(_310_)
);

OAI21X1 _855_ (
    .A(_161__bF$buf7),
    .B(_310_),
    .C(_589_[8]),
    .Y(_311_)
);

OAI21X1 _856_ (
    .A(_158_),
    .B(_309_),
    .C(_311_),
    .Y(_42_)
);

OAI21X1 _857_ (
    .A(_161__bF$buf6),
    .B(_310_),
    .C(_589_[9]),
    .Y(_312_)
);

OAI21X1 _858_ (
    .A(_176_),
    .B(_309_),
    .C(_312_),
    .Y(_43_)
);

OAI21X1 _859_ (
    .A(_161__bF$buf5),
    .B(_310_),
    .C(_589_[10]),
    .Y(_313_)
);

OAI21X1 _860_ (
    .A(_190_),
    .B(_309_),
    .C(_313_),
    .Y(_44_)
);

OAI21X1 _861_ (
    .A(_161__bF$buf4),
    .B(_310_),
    .C(_589_[11]),
    .Y(_314_)
);

OAI21X1 _862_ (
    .A(_204_),
    .B(_309_),
    .C(_314_),
    .Y(_45_)
);

OAI21X1 _863_ (
    .A(_161__bF$buf3),
    .B(_310_),
    .C(_589_[12]),
    .Y(_315_)
);

OAI21X1 _864_ (
    .A(_218_),
    .B(_309_),
    .C(_315_),
    .Y(_46_)
);

OAI21X1 _865_ (
    .A(_161__bF$buf2),
    .B(_310_),
    .C(_589_[13]),
    .Y(_316_)
);

OAI21X1 _866_ (
    .A(_232_),
    .B(_309_),
    .C(_316_),
    .Y(_47_)
);

OAI21X1 _867_ (
    .A(_161__bF$buf1),
    .B(_310_),
    .C(_589_[14]),
    .Y(_317_)
);

OAI21X1 _868_ (
    .A(_245_),
    .B(_309_),
    .C(_317_),
    .Y(_48_)
);

OAI21X1 _869_ (
    .A(_161__bF$buf0),
    .B(_310_),
    .C(_589_[15]),
    .Y(_318_)
);

OAI21X1 _870_ (
    .A(_257_),
    .B(_309_),
    .C(_318_),
    .Y(_49_)
);

NOR2X1 _871_ (
    .A(_307_),
    .B(_125_),
    .Y(_319_)
);

OAI21X1 _872_ (
    .A(_120_),
    .B(_123_),
    .C(_319_),
    .Y(_320_)
);

INVX4 _873_ (
    .A(_319_),
    .Y(_321_)
);

OAI21X1 _874_ (
    .A(_161__bF$buf7),
    .B(_321_),
    .C(_589_[16]),
    .Y(_322_)
);

OAI21X1 _875_ (
    .A(_158_),
    .B(_320_),
    .C(_322_),
    .Y(_50_)
);

OAI21X1 _876_ (
    .A(_161__bF$buf6),
    .B(_321_),
    .C(_589_[17]),
    .Y(_323_)
);

OAI21X1 _877_ (
    .A(_176_),
    .B(_320_),
    .C(_323_),
    .Y(_51_)
);

OAI21X1 _878_ (
    .A(_161__bF$buf5),
    .B(_321_),
    .C(_589_[18]),
    .Y(_324_)
);

OAI21X1 _879_ (
    .A(_190_),
    .B(_320_),
    .C(_324_),
    .Y(_52_)
);

OAI21X1 _880_ (
    .A(_161__bF$buf4),
    .B(_321_),
    .C(_589_[19]),
    .Y(_325_)
);

OAI21X1 _881_ (
    .A(_204_),
    .B(_320_),
    .C(_325_),
    .Y(_53_)
);

OAI21X1 _882_ (
    .A(_161__bF$buf3),
    .B(_321_),
    .C(_589_[20]),
    .Y(_326_)
);

OAI21X1 _883_ (
    .A(_218_),
    .B(_320_),
    .C(_326_),
    .Y(_54_)
);

OAI21X1 _884_ (
    .A(_161__bF$buf2),
    .B(_321_),
    .C(_589_[21]),
    .Y(_327_)
);

OAI21X1 _885_ (
    .A(_232_),
    .B(_320_),
    .C(_327_),
    .Y(_55_)
);

OAI21X1 _886_ (
    .A(_161__bF$buf1),
    .B(_321_),
    .C(_589_[22]),
    .Y(_328_)
);

OAI21X1 _887_ (
    .A(_245_),
    .B(_320_),
    .C(_328_),
    .Y(_56_)
);

OAI21X1 _888_ (
    .A(_161__bF$buf0),
    .B(_321_),
    .C(_589_[23]),
    .Y(_329_)
);

OAI21X1 _889_ (
    .A(_257_),
    .B(_320_),
    .C(_329_),
    .Y(_57_)
);

INVX1 _890_ (
    .A(_295_),
    .Y(_330_)
);

NAND2X1 _891_ (
    .A(instr[10]),
    .B(_330_),
    .Y(_331_)
);

INVX1 _892_ (
    .A(_331_),
    .Y(_332_)
);

OAI21X1 _893_ (
    .A(_120_),
    .B(_123_),
    .C(_332_),
    .Y(_333_)
);

OAI21X1 _894_ (
    .A(_161__bF$buf7),
    .B(_331_),
    .C(_590_[0]),
    .Y(_334_)
);

OAI21X1 _895_ (
    .A(_158_),
    .B(_333_),
    .C(_334_),
    .Y(_58_)
);

OAI21X1 _896_ (
    .A(_161__bF$buf6),
    .B(_331_),
    .C(_590_[1]),
    .Y(_335_)
);

OAI21X1 _897_ (
    .A(_176_),
    .B(_333_),
    .C(_335_),
    .Y(_59_)
);

OAI21X1 _898_ (
    .A(_161__bF$buf5),
    .B(_331_),
    .C(_590_[2]),
    .Y(_336_)
);

OAI21X1 _899_ (
    .A(_190_),
    .B(_333_),
    .C(_336_),
    .Y(_60_)
);

OAI21X1 _900_ (
    .A(_161__bF$buf4),
    .B(_331_),
    .C(_590_[3]),
    .Y(_337_)
);

OAI21X1 _901_ (
    .A(_204_),
    .B(_333_),
    .C(_337_),
    .Y(_61_)
);

OAI21X1 _902_ (
    .A(_161__bF$buf3),
    .B(_331_),
    .C(_590_[4]),
    .Y(_338_)
);

OAI21X1 _903_ (
    .A(_218_),
    .B(_333_),
    .C(_338_),
    .Y(_62_)
);

OAI21X1 _904_ (
    .A(_161__bF$buf2),
    .B(_331_),
    .C(_590_[5]),
    .Y(_339_)
);

OAI21X1 _905_ (
    .A(_232_),
    .B(_333_),
    .C(_339_),
    .Y(_63_)
);

OAI21X1 _906_ (
    .A(_161__bF$buf1),
    .B(_331_),
    .C(_590_[6]),
    .Y(_340_)
);

OAI21X1 _907_ (
    .A(_245_),
    .B(_333_),
    .C(_340_),
    .Y(_64_)
);

OAI21X1 _908_ (
    .A(_161__bF$buf0),
    .B(_331_),
    .C(_590_[7]),
    .Y(_341_)
);

OAI21X1 _909_ (
    .A(_257_),
    .B(_333_),
    .C(_341_),
    .Y(_65_)
);

INVX2 _910_ (
    .A(_592_[0]),
    .Y(_342_)
);

INVX1 _911_ (
    .A(instr[8]),
    .Y(_343_)
);

NAND2X1 _912_ (
    .A(\ALU_H4.cout ),
    .B(_343_),
    .Y(_344_)
);

NOR2X1 _913_ (
    .A(instr[9]),
    .B(_307_),
    .Y(_345_)
);

AOI22X1 _914_ (
    .A(_344_),
    .B(_345_),
    .C(_259_),
    .D(_152_),
    .Y(_346_)
);

NAND2X1 _915_ (
    .A(\ALU_H4.eqv ),
    .B(\ALU_L4.eqv ),
    .Y(_347_)
);

AOI22X1 _916_ (
    .A(_296_),
    .B(_347_),
    .C(_126_),
    .D(_237_),
    .Y(_348_)
);

NAND2X1 _917_ (
    .A(_346_),
    .B(_348_),
    .Y(_349_)
);

NOR2X1 _918_ (
    .A(_92_),
    .B(_97_),
    .Y(_350_)
);

NAND2X1 _919_ (
    .A(_350_),
    .B(_349_),
    .Y(_351_)
);

NOR2X1 _920_ (
    .A(_589_[0]),
    .B(_351__bF$buf0),
    .Y(_352_)
);

INVX4 _921_ (
    .A(_351__bF$buf4),
    .Y(_353_)
);

OAI21X1 _922_ (
    .A(_353_),
    .B(_342_),
    .C(_93__bF$buf4),
    .Y(_354_)
);

OAI22X1 _923_ (
    .A(_93__bF$buf3),
    .B(_342_),
    .C(_354_),
    .D(_352_),
    .Y(_66_)
);

INVX1 _924_ (
    .A(_592_[1]),
    .Y(_355_)
);

NAND2X1 _925_ (
    .A(_592_[0]),
    .B(_592_[1]),
    .Y(_356_)
);

NAND2X1 _926_ (
    .A(_342_),
    .B(_355_),
    .Y(_357_)
);

NAND3X1 _927_ (
    .A(_356_),
    .B(_357_),
    .C(_351__bF$buf3),
    .Y(_358_)
);

AOI21X1 _928_ (
    .A(_589_[1]),
    .B(_353_),
    .C(WAIT_bF$buf3),
    .Y(_359_)
);

AOI22X1 _929_ (
    .A(WAIT_bF$buf2),
    .B(_355_),
    .C(_359_),
    .D(_358_),
    .Y(_67_)
);

AND2X2 _930_ (
    .A(_592_[0]),
    .B(_592_[1]),
    .Y(_360_)
);

NAND2X1 _931_ (
    .A(_592_[2]),
    .B(_360_),
    .Y(_361_)
);

INVX1 _932_ (
    .A(_361_),
    .Y(_362_)
);

NOR2X1 _933_ (
    .A(_592_[2]),
    .B(_360_),
    .Y(_363_)
);

OAI21X1 _934_ (
    .A(_362_),
    .B(_363_),
    .C(_351__bF$buf2),
    .Y(_364_)
);

OAI21X1 _935_ (
    .A(_589_[2]),
    .B(_351__bF$buf1),
    .C(_364_),
    .Y(_365_)
);

NAND2X1 _936_ (
    .A(WAIT_bF$buf1),
    .B(_592_[2]),
    .Y(_366_)
);

OAI21X1 _937_ (
    .A(_365_),
    .B(WAIT_bF$buf0),
    .C(_366_),
    .Y(_68_)
);

NAND2X1 _938_ (
    .A(_592_[2]),
    .B(_592_[3]),
    .Y(_367_)
);

NOR2X1 _939_ (
    .A(_356_),
    .B(_367_),
    .Y(_368_)
);

NOR2X1 _940_ (
    .A(_592_[3]),
    .B(_362_),
    .Y(_369_)
);

OAI21X1 _941_ (
    .A(_368_),
    .B(_369_),
    .C(_351__bF$buf0),
    .Y(_370_)
);

OAI21X1 _942_ (
    .A(_589_[3]),
    .B(_351__bF$buf4),
    .C(_370_),
    .Y(_371_)
);

NAND2X1 _943_ (
    .A(WAIT_bF$buf4),
    .B(_592_[3]),
    .Y(_372_)
);

OAI21X1 _944_ (
    .A(_371_),
    .B(WAIT_bF$buf3),
    .C(_372_),
    .Y(_69_)
);

NAND2X1 _945_ (
    .A(WAIT_bF$buf2),
    .B(_592_[4]),
    .Y(_373_)
);

XOR2X1 _946_ (
    .A(_368_),
    .B(_592_[4]),
    .Y(_374_)
);

MUX2X1 _947_ (
    .A(_374_),
    .B(_589_[4]),
    .S(_351__bF$buf3),
    .Y(_375_)
);

OAI21X1 _948_ (
    .A(_375_),
    .B(WAIT_bF$buf1),
    .C(_373_),
    .Y(_70_)
);

AND2X2 _949_ (
    .A(_592_[2]),
    .B(_592_[3]),
    .Y(_376_)
);

AND2X2 _950_ (
    .A(_592_[4]),
    .B(_592_[5]),
    .Y(_377_)
);

NAND3X1 _951_ (
    .A(_360_),
    .B(_376_),
    .C(_377_),
    .Y(_378_)
);

INVX1 _952_ (
    .A(_378_),
    .Y(_379_)
);

AOI21X1 _953_ (
    .A(_592_[4]),
    .B(_368_),
    .C(_592_[5]),
    .Y(_380_)
);

OAI21X1 _954_ (
    .A(_379_),
    .B(_380_),
    .C(_351__bF$buf2),
    .Y(_381_)
);

OAI21X1 _955_ (
    .A(_589_[5]),
    .B(_351__bF$buf1),
    .C(_381_),
    .Y(_382_)
);

NAND2X1 _956_ (
    .A(WAIT_bF$buf0),
    .B(_592_[5]),
    .Y(_383_)
);

OAI21X1 _957_ (
    .A(_382_),
    .B(WAIT_bF$buf4),
    .C(_383_),
    .Y(_71_)
);

NAND2X1 _958_ (
    .A(WAIT_bF$buf3),
    .B(_592_[6]),
    .Y(_384_)
);

XNOR2X1 _959_ (
    .A(_378_),
    .B(_592_[6]),
    .Y(_385_)
);

MUX2X1 _960_ (
    .A(_385_),
    .B(_589_[6]),
    .S(_351__bF$buf0),
    .Y(_386_)
);

OAI21X1 _961_ (
    .A(_386_),
    .B(WAIT_bF$buf2),
    .C(_384_),
    .Y(_72_)
);

NAND2X1 _962_ (
    .A(WAIT_bF$buf1),
    .B(_592_[7]),
    .Y(_387_)
);

INVX1 _963_ (
    .A(_97_),
    .Y(_388_)
);

NAND3X1 _964_ (
    .A(_102_),
    .B(_388_),
    .C(_349_),
    .Y(_389_)
);

NAND2X1 _965_ (
    .A(_592_[6]),
    .B(_379_),
    .Y(_390_)
);

XOR2X1 _966_ (
    .A(_390_),
    .B(_592_[7]),
    .Y(_391_)
);

NAND2X1 _967_ (
    .A(_351__bF$buf4),
    .B(_391_),
    .Y(_392_)
);

OAI21X1 _968_ (
    .A(_589_[7]),
    .B(_389_),
    .C(_392_),
    .Y(_393_)
);

OAI21X1 _969_ (
    .A(_393_),
    .B(WAIT_bF$buf0),
    .C(_387_),
    .Y(_73_)
);

NAND2X1 _970_ (
    .A(_592_[6]),
    .B(_592_[7]),
    .Y(_394_)
);

NOR2X1 _971_ (
    .A(_394_),
    .B(_378_),
    .Y(_395_)
);

NOR2X1 _972_ (
    .A(_592_[8]),
    .B(_395_),
    .Y(_396_)
);

INVX1 _973_ (
    .A(_592_[8]),
    .Y(_397_)
);

NAND2X1 _974_ (
    .A(_592_[4]),
    .B(_592_[5]),
    .Y(_398_)
);

NOR2X1 _975_ (
    .A(_367_),
    .B(_398_),
    .Y(_399_)
);

NOR2X1 _976_ (
    .A(_356_),
    .B(_394_),
    .Y(_400_)
);

NAND2X1 _977_ (
    .A(_399_),
    .B(_400_),
    .Y(_401_)
);

NOR2X1 _978_ (
    .A(_397_),
    .B(_401_),
    .Y(_402_)
);

OAI21X1 _979_ (
    .A(_396_),
    .B(_402_),
    .C(_351__bF$buf3),
    .Y(_403_)
);

OAI21X1 _980_ (
    .A(_589_[8]),
    .B(_351__bF$buf2),
    .C(_403_),
    .Y(_404_)
);

NAND2X1 _981_ (
    .A(WAIT_bF$buf4),
    .B(_592_[8]),
    .Y(_405_)
);

OAI21X1 _982_ (
    .A(_404_),
    .B(WAIT_bF$buf3),
    .C(_405_),
    .Y(_74_)
);

INVX1 _983_ (
    .A(_394_),
    .Y(_406_)
);

NAND3X1 _984_ (
    .A(_377_),
    .B(_406_),
    .C(_368_),
    .Y(_407_)
);

NAND2X1 _985_ (
    .A(_592_[8]),
    .B(_592_[9]),
    .Y(_408_)
);

NOR2X1 _986_ (
    .A(_408_),
    .B(_407_),
    .Y(_409_)
);

AOI21X1 _987_ (
    .A(_592_[8]),
    .B(_395_),
    .C(_592_[9]),
    .Y(_410_)
);

OAI21X1 _988_ (
    .A(_409_),
    .B(_410_),
    .C(_351__bF$buf1),
    .Y(_411_)
);

OAI21X1 _989_ (
    .A(_589_[9]),
    .B(_351__bF$buf0),
    .C(_411_),
    .Y(_412_)
);

NAND2X1 _990_ (
    .A(WAIT_bF$buf2),
    .B(_592_[9]),
    .Y(_413_)
);

OAI21X1 _991_ (
    .A(_412_),
    .B(WAIT_bF$buf1),
    .C(_413_),
    .Y(_75_)
);

INVX1 _992_ (
    .A(_592_[10]),
    .Y(_414_)
);

OAI21X1 _993_ (
    .A(_407_),
    .B(_408_),
    .C(_414_),
    .Y(_415_)
);

NAND2X1 _994_ (
    .A(_592_[10]),
    .B(_409_),
    .Y(_416_)
);

AOI21X1 _995_ (
    .A(_415_),
    .B(_416_),
    .C(_353_),
    .Y(_417_)
);

OAI21X1 _996_ (
    .A(_351__bF$buf4),
    .B(_589_[10]),
    .C(_93__bF$buf2),
    .Y(_418_)
);

OAI22X1 _997_ (
    .A(_93__bF$buf1),
    .B(_414_),
    .C(_417_),
    .D(_418_),
    .Y(_76_)
);

NAND2X1 _998_ (
    .A(WAIT_bF$buf0),
    .B(_592_[11]),
    .Y(_419_)
);

NOR2X1 _999_ (
    .A(_398_),
    .B(_394_),
    .Y(_420_)
);

endmodule
