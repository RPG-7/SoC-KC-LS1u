//配备FSB8的“最小化”KC-LS1u应用处理器
//i8088风格
//目标器件GW1N-1
module MIN_LS1u
(

);




endmodule 