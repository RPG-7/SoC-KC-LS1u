`define VENDOR_ANLOGIC
