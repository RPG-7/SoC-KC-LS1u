`define VENDOR_ASIC