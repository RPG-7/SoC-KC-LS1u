`define VENDOR_GOWIN
