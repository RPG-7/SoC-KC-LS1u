module vga_font
(
    
);



endmodule