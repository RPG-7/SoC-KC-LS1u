`define VENDOR_SIMU