`define VENDOR_ALTERA
