module SoC_LS1u
(
    input clk,
    input rst,
    output qsel,
    inout [3:0]qspi,
    inout [2:0]gpio,
    output [3:0]spi_devsel,
    output spi_cs,
    output mosi,
    output mclk,
    input miso

);


endmodule
