module SoC_LS1u
(
    
);


endmodule
